module neorv32_cpu_cp_muldiv_32_3f29546453678b855931c174a97d6c0894b8f546
  (input  clk_i,
   input  rstn_i,
   input  ctrl_i_rf_wb_en,
   input  [4:0] ctrl_i_rf_rs1,
   input  [4:0] ctrl_i_rf_rs2,
   input  [4:0] ctrl_i_rf_rs3,
   input  [4:0] ctrl_i_rf_rd,
   input  [1:0] ctrl_i_rf_mux,
   input  ctrl_i_rf_zero_we,
   input  [2:0] ctrl_i_alu_op,
   input  ctrl_i_alu_opa_mux,
   input  ctrl_i_alu_opb_mux,
   input  ctrl_i_alu_unsigned,
   input  [2:0] ctrl_i_alu_frm,
   input  [5:0] ctrl_i_alu_cp_trig,
   input  ctrl_i_bus_req,
   input  ctrl_i_bus_mo_we,
   input  ctrl_i_bus_fence,
   input  ctrl_i_bus_fencei,
   input  ctrl_i_bus_priv,
   input  [2:0] ctrl_i_ir_funct3,
   input  [11:0] ctrl_i_ir_funct12,
   input  [6:0] ctrl_i_ir_opcode,
   input  ctrl_i_cpu_priv,
   input  ctrl_i_cpu_sleep,
   input  ctrl_i_cpu_trap,
   input  ctrl_i_cpu_debug,
   input  start_i,
   input  [31:0] rs1_i,
   input  [31:0] rs2_i,
   output [31:0] res_o,
   output valid_o);
  wire [69:0] n12302_o;
  wire [48:0] ctrl;
  wire [162:0] div;
  wire [230:0] mul;
  wire n12306_o;
  wire [1:0] n12315_o;
  wire [2:0] n12316_o;
  wire [1:0] n12319_o;
  wire n12321_o;
  wire n12322_o;
  wire n12323_o;
  wire n12324_o;
  wire n12331_o;
  wire n12333_o;
  wire n12335_o;
  wire n12336_o;
  wire n12337_o;
  wire n12338_o;
  wire n12339_o;
  wire n12340_o;
  wire n12341_o;
  wire n12342_o;
  wire n12343_o;
  wire n12344_o;
  wire n12345_o;
  wire n12346_o;
  wire n12347_o;
  wire n12348_o;
  wire n12349_o;
  wire n12350_o;
  wire n12351_o;
  wire n12352_o;
  wire n12353_o;
  wire n12354_o;
  wire n12355_o;
  wire n12356_o;
  wire n12357_o;
  wire n12358_o;
  wire n12359_o;
  wire n12360_o;
  wire n12361_o;
  wire n12362_o;
  wire n12363_o;
  wire n12364_o;
  wire n12365_o;
  wire n12366_o;
  wire n12367_o;
  wire n12368_o;
  wire n12369_o;
  wire n12370_o;
  wire n12371_o;
  wire n12372_o;
  wire n12373_o;
  wire n12374_o;
  wire n12375_o;
  wire n12376_o;
  wire n12377_o;
  wire n12378_o;
  wire n12379_o;
  wire n12380_o;
  wire n12381_o;
  wire n12382_o;
  wire n12383_o;
  wire n12384_o;
  wire n12385_o;
  wire n12386_o;
  wire n12387_o;
  wire n12388_o;
  wire n12389_o;
  wire n12390_o;
  wire n12391_o;
  wire n12392_o;
  wire n12393_o;
  wire n12394_o;
  wire n12395_o;
  wire n12396_o;
  wire n12397_o;
  wire [1:0] n12398_o;
  wire n12400_o;
  wire n12401_o;
  wire n12403_o;
  wire n12404_o;
  wire n12405_o;
  wire n12406_o;
  wire n12407_o;
  wire [31:0] n12409_o;
  wire [31:0] n12410_o;
  wire [1:0] n12414_o;
  wire [1:0] n12415_o;
  wire [31:0] n12416_o;
  wire [31:0] n12417_o;
  wire n12418_o;
  wire n12419_o;
  wire n12421_o;
  wire [4:0] n12422_o;
  wire [4:0] n12424_o;
  wire [4:0] n12426_o;
  wire n12432_o;
  wire n12434_o;
  wire n12436_o;
  wire n12437_o;
  wire n12438_o;
  wire n12439_o;
  wire n12440_o;
  wire n12441_o;
  wire n12442_o;
  wire n12443_o;
  wire n12444_o;
  wire n12445_o;
  wire n12446_o;
  wire [1:0] n12448_o;
  wire [1:0] n12449_o;
  wire n12451_o;
  wire n12455_o;
  wire [2:0] n12457_o;
  reg [1:0] n12458_o;
  wire [4:0] n12459_o;
  reg [4:0] n12460_o;
  wire [2:0] n12461_o;
  reg [2:0] n12462_o;
  reg n12463_o;
  wire [31:0] n12464_o;
  reg [31:0] n12465_o;
  wire n12466_o;
  reg n12467_o;
  wire [6:0] n12468_o;
  wire [32:0] n12469_o;
  wire [6:0] n12478_o;
  wire [32:0] n12479_o;
  wire [1:0] n12486_o;
  wire n12488_o;
  wire n12489_o;
  wire [2:0] n12491_o;
  wire n12493_o;
  wire n12494_o;
  wire [2:0] n12497_o;
  wire n12499_o;
  wire [2:0] n12500_o;
  wire n12502_o;
  wire n12503_o;
  wire [2:0] n12504_o;
  wire n12506_o;
  wire n12507_o;
  wire [2:0] n12508_o;
  wire n12510_o;
  wire n12511_o;
  wire n12512_o;
  wire [2:0] n12515_o;
  wire n12517_o;
  wire [2:0] n12518_o;
  wire n12520_o;
  wire n12521_o;
  wire [2:0] n12522_o;
  wire n12524_o;
  wire n12525_o;
  wire n12526_o;
  wire n12529_o;
  wire n12530_o;
  wire n12531_o;
  wire n12532_o;
  wire n12535_o;
  wire n12536_o;
  wire n12537_o;
  wire n12544_o;
  wire [1:0] n12546_o;
  wire n12548_o;
  wire [1:0] n12549_o;
  wire n12551_o;
  wire n12552_o;
  wire [32:0] n12553_o;
  wire [30:0] n12554_o;
  wire [63:0] n12555_o;
  wire [63:0] n12556_o;
  wire [63:0] n12557_o;
  wire [63:0] n12558_o;
  wire [63:0] n12559_o;
  wire n12564_o;
  wire [1:0] n12565_o;
  wire n12567_o;
  wire n12568_o;
  wire n12569_o;
  wire n12570_o;
  wire [31:0] n12571_o;
  wire [32:0] n12572_o;
  wire n12573_o;
  wire n12574_o;
  wire n12575_o;
  wire [32:0] n12576_o;
  wire [32:0] n12577_o;
  wire n12578_o;
  wire [31:0] n12579_o;
  wire [32:0] n12580_o;
  wire n12581_o;
  wire n12582_o;
  wire n12583_o;
  wire [32:0] n12584_o;
  wire [32:0] n12585_o;
  wire [32:0] n12586_o;
  wire n12587_o;
  wire [31:0] n12588_o;
  wire [32:0] n12589_o;
  wire [32:0] n12590_o;
  wire n12592_o;
  wire n12593_o;
  wire n12594_o;
  wire n12597_o;
  wire n12598_o;
  wire n12599_o;
  wire n12600_o;
  wire [31:0] n12602_o;
  wire [31:0] n12603_o;
  wire [1:0] n12605_o;
  wire n12607_o;
  wire [1:0] n12608_o;
  wire n12610_o;
  wire n12611_o;
  wire [30:0] n12612_o;
  wire n12613_o;
  wire n12614_o;
  wire [31:0] n12615_o;
  wire n12616_o;
  wire n12617_o;
  wire [31:0] n12618_o;
  wire [30:0] n12619_o;
  wire n12620_o;
  wire [31:0] n12621_o;
  wire [31:0] n12622_o;
  wire [63:0] n12623_o;
  wire [63:0] n12624_o;
  wire [63:0] n12625_o;
  wire [63:0] n12626_o;
  wire [63:0] n12627_o;
  wire [30:0] n12631_o;
  wire [31:0] n12633_o;
  wire n12634_o;
  wire [32:0] n12635_o;
  wire [31:0] n12636_o;
  wire [32:0] n12638_o;
  wire [32:0] n12639_o;
  wire [31:0] n12640_o;
  wire [2:0] n12641_o;
  wire n12643_o;
  wire [2:0] n12644_o;
  wire n12646_o;
  wire n12647_o;
  wire [31:0] n12648_o;
  wire [31:0] n12649_o;
  wire [31:0] n12650_o;
  wire [31:0] n12652_o;
  wire n12653_o;
  wire [31:0] n12654_o;
  wire [31:0] n12655_o;
  wire n12657_o;
  wire [2:0] n12658_o;
  wire [31:0] n12659_o;
  wire n12661_o;
  wire [31:0] n12662_o;
  wire n12664_o;
  wire n12666_o;
  wire n12667_o;
  wire n12669_o;
  wire n12670_o;
  wire [31:0] n12671_o;
  wire [1:0] n12672_o;
  reg [31:0] n12673_o;
  wire [31:0] n12675_o;
  reg [32:0] n12678_q;
  reg [2:0] n12679_q;
  reg [6:0] n12680_q;
  wire [48:0] n12681_o;
  reg [63:0] n12682_q;
  reg n12683_q;
  wire [162:0] n12684_o;
  reg [63:0] n12685_q;
  wire [230:0] n12686_o;
  assign res_o = n12675_o;
  assign valid_o = n12489_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:60:5  */
  assign n12302_o = {ctrl_i_cpu_debug, ctrl_i_cpu_trap, ctrl_i_cpu_sleep, ctrl_i_cpu_priv, ctrl_i_ir_opcode, ctrl_i_ir_funct12, ctrl_i_ir_funct3, ctrl_i_bus_priv, ctrl_i_bus_fencei, ctrl_i_bus_fence, ctrl_i_bus_mo_we, ctrl_i_bus_req, ctrl_i_alu_cp_trig, ctrl_i_alu_frm, ctrl_i_alu_unsigned, ctrl_i_alu_opb_mux, ctrl_i_alu_opa_mux, ctrl_i_alu_op, ctrl_i_rf_zero_we, ctrl_i_rf_mux, ctrl_i_rf_rd, ctrl_i_rf_rs3, ctrl_i_rf_rs2, ctrl_i_rf_rs1, ctrl_i_rf_wb_en};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:92:10  */
  assign ctrl = n12681_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:104:10  */
  assign div = n12684_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:116:10  */
  assign mul = n12686_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:124:16  */
  assign n12306_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:136:17  */
  assign n12315_o = ctrl[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:140:33  */
  assign n12316_o = ctrl[9:7];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:145:29  */
  assign n12319_o = ctrl[8:7];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:145:42  */
  assign n12321_o = n12319_o == 2'b00;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:146:39  */
  assign n12322_o = rs1_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:146:61  */
  assign n12323_o = rs2_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:146:52  */
  assign n12324_o = n12322_o ^ n12323_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12331_o = rs2_i[31];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12333_o = 1'b0 | n12331_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12335_o = rs2_i[30];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12336_o = n12333_o | n12335_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12337_o = rs2_i[29];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12338_o = n12336_o | n12337_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12339_o = rs2_i[28];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12340_o = n12338_o | n12339_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12341_o = rs2_i[27];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12342_o = n12340_o | n12341_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12343_o = rs2_i[26];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12344_o = n12342_o | n12343_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12345_o = rs2_i[25];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12346_o = n12344_o | n12345_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12347_o = rs2_i[24];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12348_o = n12346_o | n12347_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12349_o = rs2_i[23];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12350_o = n12348_o | n12349_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12351_o = rs2_i[22];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12352_o = n12350_o | n12351_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12353_o = rs2_i[21];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12354_o = n12352_o | n12353_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12355_o = rs2_i[20];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12356_o = n12354_o | n12355_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12357_o = rs2_i[19];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12358_o = n12356_o | n12357_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12359_o = rs2_i[18];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12360_o = n12358_o | n12359_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12361_o = rs2_i[17];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12362_o = n12360_o | n12361_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12363_o = rs2_i[16];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12364_o = n12362_o | n12363_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12365_o = rs2_i[15];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12366_o = n12364_o | n12365_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12367_o = rs2_i[14];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12368_o = n12366_o | n12367_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12369_o = rs2_i[13];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12370_o = n12368_o | n12369_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12371_o = rs2_i[12];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12372_o = n12370_o | n12371_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12373_o = rs2_i[11];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12374_o = n12372_o | n12373_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12375_o = rs2_i[10];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12376_o = n12374_o | n12375_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12377_o = rs2_i[9];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12378_o = n12376_o | n12377_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12379_o = rs2_i[8];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12380_o = n12378_o | n12379_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12381_o = rs2_i[7];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12382_o = n12380_o | n12381_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12383_o = rs2_i[6];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12384_o = n12382_o | n12383_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12385_o = rs2_i[5];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12386_o = n12384_o | n12385_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12387_o = rs2_i[4];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12388_o = n12386_o | n12387_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12389_o = rs2_i[3];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12390_o = n12388_o | n12389_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12391_o = rs2_i[2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12392_o = n12390_o | n12391_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12393_o = rs2_i[1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12394_o = n12392_o | n12393_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12395_o = rs2_i[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12396_o = n12394_o | n12395_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:146:75  */
  assign n12397_o = n12324_o & n12396_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:147:32  */
  assign n12398_o = ctrl[8:7];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:147:45  */
  assign n12400_o = n12398_o == 2'b10;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:148:38  */
  assign n12401_o = rs1_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:147:15  */
  assign n12403_o = n12400_o ? n12401_o : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:145:15  */
  assign n12404_o = n12321_o ? n12397_o : n12403_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:153:25  */
  assign n12405_o = rs2_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:153:47  */
  assign n12406_o = ctrl[15];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:153:38  */
  assign n12407_o = n12405_o & n12406_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:154:53  */
  assign n12409_o = 32'b00000000000000000000000000000000 - rs2_i;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:153:15  */
  assign n12410_o = n12407_o ? n12409_o : rs2_i;
  assign n12414_o = ctrl[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:142:11  */
  assign n12415_o = start_i ? 2'b01 : n12414_o;
  assign n12416_o = ctrl[48:17];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:142:11  */
  assign n12417_o = start_i ? n12410_o : n12416_o;
  assign n12418_o = div[1];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:142:11  */
  assign n12419_o = start_i ? n12404_o : n12418_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:138:9  */
  assign n12421_o = n12315_o == 2'b00;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:168:55  */
  assign n12422_o = ctrl[6:2];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:168:60  */
  assign n12424_o = n12422_o - 5'b00001;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:169:32  */
  assign n12426_o = ctrl[6:2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12432_o = n12426_o[4];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12434_o = 1'b0 | n12432_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12436_o = n12426_o[3];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12437_o = n12434_o | n12436_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12438_o = n12426_o[2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12439_o = n12437_o | n12438_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12440_o = n12426_o[1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12441_o = n12439_o | n12440_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12442_o = n12426_o[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12443_o = n12441_o | n12442_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:169:37  */
  assign n12444_o = ~n12443_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:169:55  */
  assign n12445_o = n12302_o[68];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:169:44  */
  assign n12446_o = n12444_o | n12445_o;
  assign n12448_o = ctrl[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:169:11  */
  assign n12449_o = n12446_o ? 2'b10 : n12448_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:167:9  */
  assign n12451_o = n12315_o == 2'b01;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:173:9  */
  assign n12455_o = n12315_o == 2'b10;
  assign n12457_o = {n12455_o, n12451_o, n12421_o};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:136:7  */
  always @*
    case (n12457_o)
      3'b100: n12458_o = 2'b00;
      3'b010: n12458_o = n12449_o;
      3'b001: n12458_o = n12415_o;
      default: n12458_o = 2'b00;
    endcase
  assign n12459_o = ctrl[6:2];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:136:7  */
  always @*
    case (n12457_o)
      3'b100: n12460_o = n12459_o;
      3'b010: n12460_o = n12424_o;
      3'b001: n12460_o = 5'b11110;
      default: n12460_o = n12459_o;
    endcase
  assign n12461_o = ctrl[12:10];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:136:7  */
  always @*
    case (n12457_o)
      3'b100: n12462_o = n12461_o;
      3'b010: n12462_o = n12461_o;
      3'b001: n12462_o = n12316_o;
      default: n12462_o = n12461_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:136:7  */
  always @*
    case (n12457_o)
      3'b100: n12463_o = 1'b1;
      3'b010: n12463_o = 1'b0;
      3'b001: n12463_o = 1'b0;
      default: n12463_o = 1'b0;
    endcase
  assign n12464_o = ctrl[48:17];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:136:7  */
  always @*
    case (n12457_o)
      3'b100: n12465_o = n12464_o;
      3'b010: n12465_o = n12464_o;
      3'b001: n12465_o = n12417_o;
      default: n12465_o = n12464_o;
    endcase
  assign n12466_o = div[1];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:136:7  */
  always @*
    case (n12457_o)
      3'b100: n12467_o = n12466_o;
      3'b010: n12467_o = n12466_o;
      3'b001: n12467_o = n12419_o;
      default: n12467_o = n12466_o;
    endcase
  assign n12468_o = {n12460_o, n12458_o};
  assign n12469_o = {n12465_o, n12463_o};
  assign n12478_o = {5'b00000, 2'b00};
  assign n12479_o = {32'b00000000000000000000000000000000, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:184:29  */
  assign n12486_o = ctrl[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:184:35  */
  assign n12488_o = n12486_o == 2'b10;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:184:18  */
  assign n12489_o = n12488_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:187:24  */
  assign n12491_o = n12302_o[46:44];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:188:43  */
  assign n12493_o = n12302_o[46];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:188:21  */
  assign n12494_o = n12493_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:191:40  */
  assign n12497_o = ctrl[9:7];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:191:46  */
  assign n12499_o = n12497_o == 3'b001;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:191:71  */
  assign n12500_o = ctrl[9:7];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:191:77  */
  assign n12502_o = n12500_o == 3'b010;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:191:62  */
  assign n12503_o = n12499_o | n12502_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:192:40  */
  assign n12504_o = ctrl[9:7];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:192:46  */
  assign n12506_o = n12504_o == 3'b100;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:191:95  */
  assign n12507_o = n12503_o | n12506_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:192:70  */
  assign n12508_o = ctrl[9:7];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:192:76  */
  assign n12510_o = n12508_o == 3'b110;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:192:61  */
  assign n12511_o = n12507_o | n12510_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:191:29  */
  assign n12512_o = n12511_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:193:40  */
  assign n12515_o = ctrl[9:7];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:193:46  */
  assign n12517_o = n12515_o == 3'b001;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:194:40  */
  assign n12518_o = ctrl[9:7];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:194:46  */
  assign n12520_o = n12518_o == 3'b100;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:193:62  */
  assign n12521_o = n12517_o | n12520_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:194:70  */
  assign n12522_o = ctrl[9:7];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:194:76  */
  assign n12524_o = n12522_o == 3'b110;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:194:61  */
  assign n12525_o = n12521_o | n12524_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:193:29  */
  assign n12526_o = n12525_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:197:51  */
  assign n12529_o = ctrl[13];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:197:54  */
  assign n12530_o = ~n12529_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:197:41  */
  assign n12531_o = start_i & n12530_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:197:20  */
  assign n12532_o = n12531_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:198:51  */
  assign n12535_o = ctrl[13];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:198:41  */
  assign n12536_o = start_i & n12535_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:198:20  */
  assign n12537_o = n12536_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:241:17  */
  assign n12544_o = mul[0];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:244:21  */
  assign n12546_o = ctrl[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:244:27  */
  assign n12548_o = n12546_o == 2'b01;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:244:46  */
  assign n12549_o = ctrl[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:244:52  */
  assign n12551_o = n12549_o == 2'b10;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:244:37  */
  assign n12552_o = n12548_o | n12551_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:245:44  */
  assign n12553_o = mul[97:65];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:246:45  */
  assign n12554_o = mul[32:2];
  assign n12555_o = {n12553_o, n12554_o};
  assign n12556_o = mul[64:1];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:244:9  */
  assign n12557_o = n12552_o ? n12555_o : n12556_o;
  assign n12558_o = {32'b00000000000000000000000000000000, rs1_i};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:241:9  */
  assign n12559_o = n12544_o ? n12558_o : n12557_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:254:19  */
  assign n12564_o = mul[1];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:255:18  */
  assign n12565_o = ctrl[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:255:24  */
  assign n12567_o = n12565_o == 2'b10;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:255:44  */
  assign n12568_o = ctrl[14];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:255:34  */
  assign n12569_o = n12567_o & n12568_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:256:53  */
  assign n12570_o = mul[98];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:256:70  */
  assign n12571_o = mul[64:33];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:256:60  */
  assign n12572_o = {n12570_o, n12571_o};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:256:103  */
  assign n12573_o = rs2_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:256:125  */
  assign n12574_o = ctrl[15];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:256:116  */
  assign n12575_o = n12573_o & n12574_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:256:140  */
  assign n12576_o = {n12575_o, rs2_i};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:256:86  */
  assign n12577_o = n12572_o - n12576_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:258:53  */
  assign n12578_o = mul[98];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:258:70  */
  assign n12579_o = mul[64:33];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:258:60  */
  assign n12580_o = {n12578_o, n12579_o};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:258:103  */
  assign n12581_o = rs2_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:258:125  */
  assign n12582_o = ctrl[15];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:258:116  */
  assign n12583_o = n12581_o & n12582_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:258:140  */
  assign n12584_o = {n12583_o, rs2_i};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:258:86  */
  assign n12585_o = n12580_o + n12584_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:255:9  */
  assign n12586_o = n12569_o ? n12577_o : n12585_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:261:24  */
  assign n12587_o = mul[98];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:261:41  */
  assign n12588_o = mul[64:33];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:261:31  */
  assign n12589_o = {n12587_o, n12588_o};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:254:7  */
  assign n12590_o = n12564_o ? n12586_o : n12589_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:266:27  */
  assign n12592_o = mul[64];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:266:52  */
  assign n12593_o = ctrl[15];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:266:43  */
  assign n12594_o = n12592_o & n12593_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:287:17  */
  assign n12597_o = div[0];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:288:21  */
  assign n12598_o = rs1_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:288:43  */
  assign n12599_o = ctrl[14];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:288:34  */
  assign n12600_o = n12598_o & n12599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:289:49  */
  assign n12602_o = 32'b00000000000000000000000000000000 - rs1_i;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:288:11  */
  assign n12603_o = n12600_o ? n12602_o : rs1_i;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:294:21  */
  assign n12605_o = ctrl[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:294:27  */
  assign n12607_o = n12605_o == 2'b01;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:294:46  */
  assign n12608_o = ctrl[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:294:52  */
  assign n12610_o = n12608_o == 2'b10;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:294:37  */
  assign n12611_o = n12607_o | n12610_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:295:39  */
  assign n12612_o = div[64:34];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:295:67  */
  assign n12613_o = div[98];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:295:56  */
  assign n12614_o = ~n12613_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:295:53  */
  assign n12615_o = {n12612_o, n12614_o};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:296:22  */
  assign n12616_o = div[98];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:296:27  */
  assign n12617_o = ~n12616_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:297:37  */
  assign n12618_o = div[97:66];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:299:43  */
  assign n12619_o = div[32:2];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:299:71  */
  assign n12620_o = div[65];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:299:57  */
  assign n12621_o = {n12619_o, n12620_o};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:296:11  */
  assign n12622_o = n12617_o ? n12618_o : n12621_o;
  assign n12623_o = {n12615_o, n12622_o};
  assign n12624_o = div[65:2];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:294:9  */
  assign n12625_o = n12611_o ? n12623_o : n12624_o;
  assign n12626_o = {n12603_o, 32'b00000000000000000000000000000000};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:287:9  */
  assign n12627_o = n12597_o ? n12626_o : n12625_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:306:62  */
  assign n12631_o = div[32:2];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:306:47  */
  assign n12633_o = {1'b0, n12631_o};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:306:90  */
  assign n12634_o = div[65];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:306:76  */
  assign n12635_o = {n12633_o, n12634_o};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:306:118  */
  assign n12636_o = ctrl[48:17];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:306:111  */
  assign n12638_o = {1'b0, n12636_o};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:306:96  */
  assign n12639_o = n12635_o - n12638_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:309:22  */
  assign n12640_o = div[65:34];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:309:42  */
  assign n12641_o = ctrl[9:7];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:309:48  */
  assign n12643_o = n12641_o == 3'b100;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:309:72  */
  assign n12644_o = ctrl[9:7];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:309:78  */
  assign n12646_o = n12644_o == 3'b101;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:309:63  */
  assign n12647_o = n12643_o | n12646_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:309:31  */
  assign n12648_o = n12647_o ? n12640_o : n12649_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:309:103  */
  assign n12649_o = div[33:2];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:310:53  */
  assign n12650_o = div[130:99];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:310:38  */
  assign n12652_o = 32'b00000000000000000000000000000000 - n12650_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:310:71  */
  assign n12653_o = div[1];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:310:61  */
  assign n12654_o = n12653_o ? n12652_o : n12655_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:310:96  */
  assign n12655_o = div[130:99];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:330:14  */
  assign n12657_o = ctrl[16];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:331:17  */
  assign n12658_o = ctrl[12:10];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:333:28  */
  assign n12659_o = mul[32:1];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:332:9  */
  assign n12661_o = n12658_o == 3'b000;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:335:28  */
  assign n12662_o = mul[64:33];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:334:9  */
  assign n12664_o = n12658_o == 3'b001;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:334:27  */
  assign n12666_o = n12658_o == 3'b010;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:334:27  */
  assign n12667_o = n12664_o | n12666_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:334:44  */
  assign n12669_o = n12658_o == 3'b011;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:334:44  */
  assign n12670_o = n12667_o | n12669_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:337:24  */
  assign n12671_o = div[162:131];
  assign n12672_o = {n12670_o, n12661_o};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:331:7  */
  always @*
    case (n12672_o)
      2'b10: n12673_o = n12662_o;
      2'b01: n12673_o = n12659_o;
      default: n12673_o = n12671_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:330:5  */
  assign n12675_o = n12657_o ? n12673_o : 32'b00000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:131:5  */
  always @(posedge clk_i or posedge n12306_o)
    if (n12306_o)
      n12678_q <= n12479_o;
    else
      n12678_q <= n12469_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:131:5  */
  always @(posedge clk_i or posedge n12306_o)
    if (n12306_o)
      n12679_q <= 3'b000;
    else
      n12679_q <= n12462_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:131:5  */
  always @(posedge clk_i or posedge n12306_o)
    if (n12306_o)
      n12680_q <= n12478_o;
    else
      n12680_q <= n12468_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:124:5  */
  assign n12681_o = {n12678_q, n12526_o, n12512_o, n12494_o, n12679_q, n12491_o, n12680_q};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:286:7  */
  always @(posedge clk_i)
    n12682_q <= n12627_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:131:5  */
  always @(posedge clk_i or posedge n12306_o)
    if (n12306_o)
      n12683_q <= 1'b0;
    else
      n12683_q <= n12467_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:124:5  */
  assign n12684_o = {n12654_o, n12648_o, n12639_o, n12682_q, n12683_q, n12537_o};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:240:7  */
  always @(posedge clk_i)
    n12685_q <= n12559_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:240:7  */
  assign n12686_o = {66'b000000000000000000000000000000000000000000000000000000000000000000, 33'b000000000000000000000000000000000, 33'b000000000000000000000000000000000, n12594_o, n12590_o, n12685_q, n12532_o};
endmodule

module neorv32_cpu_cp_shifter_32_5ba93c9db0cff93f52b521d7420e43f6eda2784f
  (input  clk_i,
   input  rstn_i,
   input  ctrl_i_rf_wb_en,
   input  [4:0] ctrl_i_rf_rs1,
   input  [4:0] ctrl_i_rf_rs2,
   input  [4:0] ctrl_i_rf_rs3,
   input  [4:0] ctrl_i_rf_rd,
   input  [1:0] ctrl_i_rf_mux,
   input  ctrl_i_rf_zero_we,
   input  [2:0] ctrl_i_alu_op,
   input  ctrl_i_alu_opa_mux,
   input  ctrl_i_alu_opb_mux,
   input  ctrl_i_alu_unsigned,
   input  [2:0] ctrl_i_alu_frm,
   input  [5:0] ctrl_i_alu_cp_trig,
   input  ctrl_i_bus_req,
   input  ctrl_i_bus_mo_we,
   input  ctrl_i_bus_fence,
   input  ctrl_i_bus_fencei,
   input  ctrl_i_bus_priv,
   input  [2:0] ctrl_i_ir_funct3,
   input  [11:0] ctrl_i_ir_funct12,
   input  [6:0] ctrl_i_ir_opcode,
   input  ctrl_i_cpu_priv,
   input  ctrl_i_cpu_sleep,
   input  ctrl_i_cpu_trap,
   input  ctrl_i_cpu_debug,
   input  start_i,
   input  [31:0] rs1_i,
   input  [4:0] shamt_i,
   output [31:0] res_o,
   output valid_o);
  wire [69:0] n12198_o;
  wire [39:0] shifter;
  wire n12202_o;
  wire n12208_o;
  wire n12210_o;
  wire n12211_o;
  wire n12212_o;
  wire n12214_o;
  wire n12215_o;
  wire n12216_o;
  wire [4:0] n12218_o;
  wire n12224_o;
  wire n12226_o;
  wire n12228_o;
  wire n12229_o;
  wire n12230_o;
  wire n12231_o;
  wire n12232_o;
  wire n12233_o;
  wire n12234_o;
  wire n12235_o;
  wire [4:0] n12236_o;
  wire [4:0] n12238_o;
  wire n12239_o;
  wire n12240_o;
  wire [30:0] n12241_o;
  wire [31:0] n12243_o;
  wire n12244_o;
  wire n12245_o;
  wire n12246_o;
  wire [30:0] n12247_o;
  wire [31:0] n12248_o;
  wire [31:0] n12249_o;
  wire [36:0] n12250_o;
  wire [36:0] n12251_o;
  wire [36:0] n12252_o;
  wire [36:0] n12253_o;
  wire [36:0] n12254_o;
  wire [1:0] n12255_o;
  wire [1:0] n12260_o;
  wire [36:0] n12261_o;
  wire [3:0] n12267_o;
  wire n12273_o;
  wire n12275_o;
  wire n12277_o;
  wire n12278_o;
  wire n12279_o;
  wire n12280_o;
  wire n12281_o;
  wire n12282_o;
  wire n12283_o;
  wire n12284_o;
  wire n12286_o;
  wire n12287_o;
  wire n12288_o;
  wire [31:0] n12289_o;
  wire n12290_o;
  wire n12291_o;
  wire n12292_o;
  wire n12293_o;
  wire [31:0] n12294_o;
  reg [36:0] n12296_q;
  reg [1:0] n12297_q;
  wire [39:0] n12298_o;
  assign res_o = n12294_o;
  assign valid_o = n12288_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:50:5  */
  assign n12198_o = {ctrl_i_cpu_debug, ctrl_i_cpu_trap, ctrl_i_cpu_sleep, ctrl_i_cpu_priv, ctrl_i_ir_opcode, ctrl_i_ir_funct12, ctrl_i_ir_funct3, ctrl_i_bus_priv, ctrl_i_bus_fencei, ctrl_i_bus_fence, ctrl_i_bus_mo_we, ctrl_i_bus_req, ctrl_i_alu_cp_trig, ctrl_i_alu_frm, ctrl_i_alu_unsigned, ctrl_i_alu_opb_mux, ctrl_i_alu_opa_mux, ctrl_i_alu_op, ctrl_i_rf_zero_we, ctrl_i_rf_mux, ctrl_i_rf_rd, ctrl_i_rf_rs3, ctrl_i_rf_rs2, ctrl_i_rf_rs1, ctrl_i_rf_wb_en};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:75:10  */
  assign shifter = n12298_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:92:18  */
  assign n12202_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:99:36  */
  assign n12208_o = shifter[0];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:102:24  */
  assign n12210_o = shifter[2];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:102:47  */
  assign n12211_o = n12198_o[68];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:102:36  */
  assign n12212_o = n12210_o | n12211_o;
  assign n12214_o = shifter[0];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:102:9  */
  assign n12215_o = n12212_o ? 1'b0 : n12214_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:100:9  */
  assign n12216_o = start_i ? 1'b1 : n12215_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:109:36  */
  assign n12218_o = shifter[7:3];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12224_o = n12218_o[4];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12226_o = 1'b0 | n12224_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12228_o = n12218_o[3];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12229_o = n12226_o | n12228_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12230_o = n12218_o[2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12231_o = n12229_o | n12230_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12232_o = n12218_o[1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12233_o = n12231_o | n12232_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12234_o = n12218_o[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12235_o = n12233_o | n12234_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:110:61  */
  assign n12236_o = shifter[7:3];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:110:66  */
  assign n12238_o = n12236_o - 5'b00001;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:111:31  */
  assign n12239_o = n12198_o[46];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:111:35  */
  assign n12240_o = ~n12239_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:112:41  */
  assign n12241_o = shifter[38:8];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:112:72  */
  assign n12243_o = {n12241_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:114:42  */
  assign n12244_o = shifter[39];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:114:83  */
  assign n12245_o = n12198_o[57];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:114:62  */
  assign n12246_o = n12244_o & n12245_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:114:103  */
  assign n12247_o = shifter[39:9];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:114:89  */
  assign n12248_o = {n12246_o, n12247_o};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:111:11  */
  assign n12249_o = n12240_o ? n12243_o : n12248_o;
  assign n12250_o = {n12249_o, n12238_o};
  assign n12251_o = shifter[39:3];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:109:9  */
  assign n12252_o = n12235_o ? n12250_o : n12251_o;
  assign n12253_o = {rs1_i, shamt_i};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:106:9  */
  assign n12254_o = start_i ? n12253_o : n12252_o;
  assign n12255_o = {n12208_o, n12216_o};
  assign n12260_o = {1'b0, 1'b0};
  assign n12261_o = {32'b00000000000000000000000000000000, 5'b00000};
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:121:54  */
  assign n12267_o = shifter[7:4];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12273_o = n12267_o[3];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12275_o = 1'b0 | n12273_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12277_o = n12267_o[2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12278_o = n12275_o | n12277_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12279_o = n12267_o[1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12280_o = n12278_o | n12279_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n12281_o = n12267_o[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n12282_o = n12280_o | n12281_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:121:83  */
  assign n12283_o = ~n12282_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:121:25  */
  assign n12284_o = n12283_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:122:29  */
  assign n12286_o = shifter[0];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:122:46  */
  assign n12287_o = shifter[2];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:122:34  */
  assign n12288_o = n12286_o & n12287_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:123:29  */
  assign n12289_o = shifter[39:8];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:123:48  */
  assign n12290_o = shifter[0];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:123:53  */
  assign n12291_o = ~n12290_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:123:73  */
  assign n12292_o = shifter[1];
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:123:60  */
  assign n12293_o = n12291_o & n12292_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:123:34  */
  assign n12294_o = n12293_o ? n12289_o : 32'b00000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:97:7  */
  always @(posedge clk_i or posedge n12202_o)
    if (n12202_o)
      n12296_q <= n12261_o;
    else
      n12296_q <= n12254_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:97:7  */
  always @(posedge clk_i or posedge n12202_o)
    if (n12202_o)
      n12297_q <= n12260_o;
    else
      n12297_q <= n12255_o;
  /* ../neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:92:7  */
  assign n12298_o = {n12296_q, n12284_o, n12297_q};
endmodule

module neorv32_cpu_decompressor_5ba93c9db0cff93f52b521d7420e43f6eda2784f
  (input  [15:0] ci_instr16_i,
   output ci_illegal_o,
   output [31:0] ci_instr32_o);
  wire n11344_o;
  wire n11345_o;
  wire n11346_o;
  wire n11347_o;
  wire n11348_o;
  wire n11349_o;
  wire n11350_o;
  wire n11351_o;
  wire n11352_o;
  wire n11353_o;
  wire n11354_o;
  wire n11355_o;
  wire n11356_o;
  wire n11357_o;
  wire n11358_o;
  wire n11359_o;
  wire n11360_o;
  wire n11361_o;
  wire n11362_o;
  wire n11363_o;
  wire n11364_o;
  wire [3:0] n11365_o;
  wire [3:0] n11366_o;
  wire [3:0] n11367_o;
  wire [3:0] n11368_o;
  wire [3:0] n11369_o;
  wire [15:0] n11370_o;
  wire [4:0] n11371_o;
  wire [20:0] n11372_o;
  wire n11375_o;
  wire n11377_o;
  wire n11379_o;
  wire n11381_o;
  wire n11383_o;
  wire n11385_o;
  wire n11387_o;
  wire n11389_o;
  wire n11391_o;
  wire n11393_o;
  wire n11395_o;
  wire [8:0] n11396_o;
  wire n11397_o;
  wire n11398_o;
  wire n11399_o;
  wire n11400_o;
  wire n11401_o;
  wire n11402_o;
  wire n11403_o;
  wire n11404_o;
  wire n11405_o;
  wire n11406_o;
  wire n11407_o;
  wire n11408_o;
  wire n11409_o;
  wire [3:0] n11410_o;
  wire [3:0] n11411_o;
  wire [3:0] n11412_o;
  wire [12:0] n11413_o;
  wire n11416_o;
  wire n11418_o;
  wire n11420_o;
  wire n11422_o;
  wire n11424_o;
  wire n11426_o;
  wire n11428_o;
  wire n11430_o;
  wire [3:0] n11431_o;
  wire [1:0] n11432_o;
  wire [2:0] n11433_o;
  localparam [1:0] n11435_o = 2'b00;
  wire n11436_o;
  wire n11437_o;
  wire n11438_o;
  wire n11439_o;
  wire n11440_o;
  localparam [4:0] n11441_o = 5'b00000;
  wire [2:0] n11443_o;
  wire [4:0] n11445_o;
  wire [2:0] n11446_o;
  wire [4:0] n11448_o;
  wire n11449_o;
  wire n11451_o;
  wire n11454_o;
  wire n11456_o;
  wire n11458_o;
  wire n11459_o;
  wire n11462_o;
  wire n11463_o;
  wire n11464_o;
  wire n11465_o;
  wire n11466_o;
  localparam [4:0] n11467_o = 5'b00000;
  wire [2:0] n11469_o;
  wire [4:0] n11471_o;
  wire [2:0] n11472_o;
  wire [4:0] n11474_o;
  wire n11475_o;
  wire n11477_o;
  wire n11480_o;
  wire n11482_o;
  wire n11484_o;
  wire n11485_o;
  wire [2:0] n11488_o;
  wire [4:0] n11490_o;
  localparam [11:0] n11492_o = 12'b000000000000;
  wire n11497_o;
  wire n11499_o;
  wire n11501_o;
  wire n11503_o;
  wire n11505_o;
  wire n11507_o;
  wire n11509_o;
  wire n11511_o;
  wire [1:0] n11512_o;
  wire [7:0] n11513_o;
  wire n11515_o;
  wire [2:0] n11516_o;
  wire n11518_o;
  wire n11519_o;
  wire [2:0] n11520_o;
  wire n11522_o;
  wire n11523_o;
  wire [2:0] n11524_o;
  wire n11526_o;
  wire n11527_o;
  wire n11530_o;
  wire [1:0] n11531_o;
  reg n11532_o;
  reg [6:0] n11533_o;
  wire [1:0] n11534_o;
  wire [1:0] n11535_o;
  reg [1:0] n11536_o;
  wire n11537_o;
  wire n11538_o;
  reg n11539_o;
  wire n11540_o;
  wire n11541_o;
  reg n11542_o;
  wire n11543_o;
  wire n11544_o;
  reg n11545_o;
  reg [2:0] n11546_o;
  reg [4:0] n11547_o;
  wire n11548_o;
  wire n11549_o;
  reg n11550_o;
  wire n11551_o;
  wire n11552_o;
  reg n11553_o;
  wire n11554_o;
  reg n11555_o;
  wire n11556_o;
  reg n11557_o;
  wire n11558_o;
  reg n11559_o;
  reg n11560_o;
  reg n11561_o;
  wire n11562_o;
  wire n11563_o;
  reg n11564_o;
  wire n11565_o;
  wire n11566_o;
  reg n11567_o;
  wire n11568_o;
  wire n11569_o;
  reg n11570_o;
  wire [1:0] n11571_o;
  wire [1:0] n11572_o;
  reg [1:0] n11573_o;
  wire n11575_o;
  wire [2:0] n11576_o;
  wire n11577_o;
  wire [4:0] n11580_o;
  wire [20:0] n11582_o;
  wire [7:0] n11583_o;
  wire [20:0] n11584_o;
  wire n11585_o;
  wire [20:0] n11586_o;
  wire [9:0] n11587_o;
  wire [20:0] n11588_o;
  wire n11589_o;
  wire n11591_o;
  wire n11593_o;
  wire n11594_o;
  wire n11595_o;
  wire n11596_o;
  wire [2:0] n11599_o;
  wire [2:0] n11601_o;
  wire [4:0] n11603_o;
  localparam [4:0] n11604_o = 5'b00000;
  wire [12:0] n11605_o;
  wire n11606_o;
  wire [12:0] n11607_o;
  wire [3:0] n11608_o;
  wire [12:0] n11609_o;
  wire [5:0] n11610_o;
  wire [12:0] n11611_o;
  wire n11612_o;
  wire n11614_o;
  wire n11616_o;
  wire n11617_o;
  wire [4:0] n11619_o;
  wire n11620_o;
  wire n11621_o;
  wire n11622_o;
  wire n11623_o;
  wire n11624_o;
  wire n11625_o;
  wire n11626_o;
  wire n11627_o;
  wire n11628_o;
  wire n11629_o;
  wire n11630_o;
  wire n11631_o;
  wire [3:0] n11632_o;
  wire [3:0] n11633_o;
  wire [3:0] n11634_o;
  wire [11:0] n11635_o;
  wire n11636_o;
  wire n11638_o;
  wire n11640_o;
  wire n11642_o;
  wire n11644_o;
  wire n11646_o;
  wire [5:0] n11647_o;
  wire n11649_o;
  wire [4:0] n11650_o;
  wire n11652_o;
  wire n11656_o;
  wire n11657_o;
  wire n11658_o;
  wire n11659_o;
  wire n11660_o;
  wire n11661_o;
  wire n11662_o;
  wire n11663_o;
  wire n11664_o;
  wire n11665_o;
  wire n11666_o;
  wire n11667_o;
  wire [3:0] n11668_o;
  wire [3:0] n11669_o;
  wire [3:0] n11670_o;
  wire [11:0] n11671_o;
  wire n11680_o;
  wire n11682_o;
  wire n11684_o;
  wire n11686_o;
  wire n11688_o;
  wire n11690_o;
  wire [1:0] n11691_o;
  wire [4:0] n11693_o;
  wire n11694_o;
  wire n11695_o;
  wire n11696_o;
  wire n11697_o;
  wire n11698_o;
  wire n11699_o;
  wire n11700_o;
  wire n11701_o;
  wire n11702_o;
  wire n11703_o;
  wire n11704_o;
  wire n11705_o;
  wire n11706_o;
  wire n11707_o;
  wire n11708_o;
  wire n11709_o;
  wire n11710_o;
  wire n11711_o;
  wire n11712_o;
  wire n11713_o;
  wire [3:0] n11714_o;
  wire [3:0] n11715_o;
  wire [3:0] n11716_o;
  wire [3:0] n11717_o;
  wire [3:0] n11718_o;
  wire [15:0] n11719_o;
  wire [19:0] n11720_o;
  wire n11721_o;
  wire n11723_o;
  wire n11725_o;
  wire n11727_o;
  wire n11729_o;
  wire n11731_o;
  wire [13:0] n11732_o;
  wire [31:0] n11733_o;
  wire [31:0] n11734_o;
  wire [31:0] n11735_o;
  wire [4:0] n11736_o;
  wire n11738_o;
  wire n11739_o;
  wire n11740_o;
  wire n11741_o;
  wire n11744_o;
  wire n11746_o;
  wire [4:0] n11747_o;
  wire [4:0] n11748_o;
  wire n11749_o;
  wire n11750_o;
  wire n11751_o;
  wire n11752_o;
  wire n11753_o;
  wire n11754_o;
  wire n11755_o;
  wire n11756_o;
  wire n11757_o;
  wire n11758_o;
  wire n11759_o;
  wire n11760_o;
  wire [3:0] n11761_o;
  wire [3:0] n11762_o;
  wire [3:0] n11763_o;
  wire [11:0] n11764_o;
  wire n11765_o;
  wire n11767_o;
  wire n11769_o;
  wire n11771_o;
  wire n11773_o;
  wire n11775_o;
  wire [5:0] n11776_o;
  wire n11778_o;
  wire [2:0] n11779_o;
  wire [4:0] n11781_o;
  wire [2:0] n11782_o;
  wire [4:0] n11784_o;
  wire [2:0] n11785_o;
  wire [4:0] n11787_o;
  wire [1:0] n11788_o;
  wire n11789_o;
  wire n11790_o;
  wire [6:0] n11793_o;
  wire n11795_o;
  wire n11796_o;
  wire n11797_o;
  wire n11798_o;
  wire n11799_o;
  wire n11800_o;
  wire n11803_o;
  wire n11805_o;
  wire n11807_o;
  wire n11808_o;
  wire n11810_o;
  wire n11811_o;
  wire n11812_o;
  wire n11813_o;
  wire n11814_o;
  wire n11815_o;
  wire n11816_o;
  wire n11817_o;
  wire n11818_o;
  wire n11819_o;
  wire n11820_o;
  wire n11821_o;
  wire [3:0] n11822_o;
  wire [3:0] n11823_o;
  wire [3:0] n11824_o;
  wire [11:0] n11825_o;
  wire n11826_o;
  wire n11828_o;
  wire n11830_o;
  wire n11832_o;
  wire n11834_o;
  wire n11836_o;
  wire [5:0] n11837_o;
  wire n11839_o;
  wire [1:0] n11841_o;
  wire n11844_o;
  wire n11848_o;
  wire n11852_o;
  wire [2:0] n11854_o;
  reg [2:0] n11855_o;
  reg [6:0] n11856_o;
  wire [1:0] n11857_o;
  reg n11859_o;
  reg [6:0] n11860_o;
  reg [2:0] n11861_o;
  wire n11862_o;
  reg n11863_o;
  wire n11864_o;
  reg n11865_o;
  wire n11866_o;
  reg n11867_o;
  wire n11868_o;
  reg n11869_o;
  wire n11870_o;
  reg n11871_o;
  wire n11872_o;
  wire n11873_o;
  reg n11874_o;
  wire [5:0] n11875_o;
  wire [5:0] n11876_o;
  reg [5:0] n11877_o;
  wire [4:0] n11882_o;
  reg n11884_o;
  wire [6:0] n11885_o;
  reg [6:0] n11886_o;
  wire n11887_o;
  wire n11888_o;
  wire n11889_o;
  wire n11890_o;
  wire n11891_o;
  reg n11892_o;
  wire [3:0] n11893_o;
  wire [3:0] n11894_o;
  wire [3:0] n11895_o;
  wire [3:0] n11896_o;
  wire [3:0] n11897_o;
  reg [3:0] n11898_o;
  wire [2:0] n11899_o;
  wire [2:0] n11900_o;
  reg [2:0] n11901_o;
  wire [4:0] n11902_o;
  wire [4:0] n11903_o;
  reg [4:0] n11904_o;
  wire n11905_o;
  wire n11906_o;
  reg n11907_o;
  wire n11908_o;
  wire n11909_o;
  wire n11910_o;
  reg n11911_o;
  wire n11912_o;
  wire n11913_o;
  wire n11914_o;
  reg n11915_o;
  wire n11916_o;
  wire n11917_o;
  wire n11918_o;
  reg n11919_o;
  wire n11920_o;
  wire n11921_o;
  wire n11922_o;
  reg n11923_o;
  wire n11924_o;
  wire n11925_o;
  wire n11926_o;
  reg n11927_o;
  wire [4:0] n11928_o;
  wire [4:0] n11929_o;
  wire [4:0] n11930_o;
  wire [4:0] n11931_o;
  wire [4:0] n11932_o;
  wire [4:0] n11933_o;
  reg [4:0] n11934_o;
  wire n11935_o;
  wire n11936_o;
  wire n11937_o;
  wire n11938_o;
  reg n11939_o;
  wire n11941_o;
  wire [2:0] n11942_o;
  wire [4:0] n11943_o;
  wire [4:0] n11944_o;
  localparam [6:0] n11946_o = 7'b0000000;
  wire n11947_o;
  wire n11948_o;
  wire n11949_o;
  wire n11950_o;
  wire n11951_o;
  wire n11952_o;
  wire n11955_o;
  wire n11957_o;
  localparam [1:0] n11958_o = 2'b00;
  wire n11959_o;
  wire n11960_o;
  wire n11961_o;
  wire n11962_o;
  wire n11963_o;
  wire n11964_o;
  wire [4:0] n11967_o;
  wire n11968_o;
  wire n11970_o;
  wire n11973_o;
  wire n11975_o;
  wire n11977_o;
  wire n11978_o;
  wire n11980_o;
  wire n11981_o;
  wire n11982_o;
  wire n11983_o;
  wire n11984_o;
  wire n11985_o;
  wire [4:0] n11988_o;
  wire n11989_o;
  wire n11991_o;
  wire n11994_o;
  wire n11996_o;
  wire n11998_o;
  wire n11999_o;
  wire n12000_o;
  wire n12001_o;
  wire [4:0] n12002_o;
  wire n12004_o;
  wire [4:0] n12006_o;
  wire [4:0] n12009_o;
  wire [4:0] n12011_o;
  wire [24:0] n12012_o;
  wire [11:0] n12013_o;
  wire [11:0] n12014_o;
  wire [11:0] n12015_o;
  wire [2:0] n12016_o;
  wire [2:0] n12018_o;
  wire [4:0] n12019_o;
  wire [4:0] n12020_o;
  wire [4:0] n12021_o;
  wire [4:0] n12023_o;
  wire [4:0] n12024_o;
  wire n12026_o;
  wire [4:0] n12027_o;
  wire n12029_o;
  wire [4:0] n12032_o;
  wire [11:0] n12034_o;
  wire [6:0] n12035_o;
  wire [6:0] n12036_o;
  wire [4:0] n12037_o;
  wire [4:0] n12039_o;
  wire [4:0] n12041_o;
  wire [11:0] n12043_o;
  wire [4:0] n12045_o;
  wire [4:0] n12046_o;
  wire [4:0] n12047_o;
  wire [24:0] n12048_o;
  wire [11:0] n12049_o;
  wire [16:0] n12050_o;
  wire [11:0] n12051_o;
  wire [11:0] n12052_o;
  wire [2:0] n12053_o;
  wire [2:0] n12055_o;
  wire [9:0] n12056_o;
  wire [9:0] n12057_o;
  wire [9:0] n12058_o;
  wire [6:0] n12059_o;
  wire [6:0] n12061_o;
  wire [31:0] n12062_o;
  wire [24:0] n12063_o;
  wire [24:0] n12064_o;
  wire [24:0] n12065_o;
  wire [6:0] n12066_o;
  wire [6:0] n12068_o;
  wire [2:0] n12069_o;
  wire n12071_o;
  wire [2:0] n12072_o;
  wire n12074_o;
  wire n12075_o;
  wire n12078_o;
  wire [2:0] n12079_o;
  reg n12080_o;
  wire [6:0] n12081_o;
  reg [6:0] n12082_o;
  wire [1:0] n12083_o;
  wire [1:0] n12084_o;
  wire [1:0] n12085_o;
  reg [1:0] n12086_o;
  wire n12087_o;
  wire n12088_o;
  wire n12089_o;
  reg n12090_o;
  wire n12091_o;
  wire n12092_o;
  wire n12093_o;
  reg n12094_o;
  wire n12095_o;
  wire n12096_o;
  wire n12097_o;
  reg n12098_o;
  wire [2:0] n12099_o;
  reg [2:0] n12100_o;
  wire [4:0] n12101_o;
  reg [4:0] n12102_o;
  wire n12103_o;
  wire n12104_o;
  wire n12105_o;
  reg n12106_o;
  wire n12107_o;
  wire n12108_o;
  wire n12109_o;
  reg n12110_o;
  wire n12111_o;
  wire n12112_o;
  reg n12113_o;
  wire n12114_o;
  wire n12115_o;
  reg n12116_o;
  wire n12117_o;
  wire n12118_o;
  reg n12119_o;
  wire n12120_o;
  wire n12121_o;
  reg n12122_o;
  wire n12123_o;
  wire n12124_o;
  reg n12125_o;
  wire n12126_o;
  wire n12127_o;
  reg n12128_o;
  wire [3:0] n12129_o;
  wire [3:0] n12130_o;
  reg [3:0] n12131_o;
  wire [1:0] n12132_o;
  reg n12133_o;
  reg [6:0] n12135_o;
  wire n12136_o;
  wire n12137_o;
  reg n12138_o;
  wire n12139_o;
  wire n12140_o;
  wire n12141_o;
  reg n12142_o;
  wire n12143_o;
  reg n12144_o;
  wire n12145_o;
  reg n12146_o;
  wire n12147_o;
  reg n12148_o;
  reg [2:0] n12149_o;
  reg [4:0] n12150_o;
  reg n12151_o;
  reg n12152_o;
  reg n12153_o;
  reg n12154_o;
  reg n12155_o;
  reg n12156_o;
  wire n12157_o;
  reg n12158_o;
  wire n12159_o;
  reg n12160_o;
  wire n12161_o;
  wire n12162_o;
  reg n12163_o;
  wire n12164_o;
  wire n12165_o;
  reg n12166_o;
  wire n12167_o;
  wire n12168_o;
  wire n12169_o;
  reg n12170_o;
  wire n12171_o;
  wire n12172_o;
  reg n12173_o;
  wire [31:0] n12197_o;
  assign ci_illegal_o = n12133_o;
  assign ci_instr32_o = n12197_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11344_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11345_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11346_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11347_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11348_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11349_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11350_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11351_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11352_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11353_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11354_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11355_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11356_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11357_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11358_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11359_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11360_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11361_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11362_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11363_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:88:39  */
  assign n11364_o = ci_instr16_i[12];
  assign n11365_o = {n11344_o, n11345_o, n11346_o, n11347_o};
  assign n11366_o = {n11348_o, n11349_o, n11350_o, n11351_o};
  assign n11367_o = {n11352_o, n11353_o, n11354_o, n11355_o};
  assign n11368_o = {n11356_o, n11357_o, n11358_o, n11359_o};
  assign n11369_o = {n11360_o, n11361_o, n11362_o, n11363_o};
  assign n11370_o = {n11365_o, n11366_o, n11367_o, n11368_o};
  assign n11371_o = {n11369_o, n11364_o};
  assign n11372_o = {n11370_o, n11371_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:90:31  */
  assign n11375_o = ci_instr16_i[3];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:91:31  */
  assign n11377_o = ci_instr16_i[4];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:92:31  */
  assign n11379_o = ci_instr16_i[5];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:93:31  */
  assign n11381_o = ci_instr16_i[11];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:94:31  */
  assign n11383_o = ci_instr16_i[2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:95:31  */
  assign n11385_o = ci_instr16_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:96:31  */
  assign n11387_o = ci_instr16_i[6];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:97:31  */
  assign n11389_o = ci_instr16_i[9];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:98:31  */
  assign n11391_o = ci_instr16_i[10];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:99:31  */
  assign n11393_o = ci_instr16_i[8];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:100:31  */
  assign n11395_o = ci_instr16_i[12];
  assign n11396_o = n11372_o[20:12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:103:39  */
  assign n11397_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:103:39  */
  assign n11398_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:103:39  */
  assign n11399_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:103:39  */
  assign n11400_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:103:39  */
  assign n11401_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:103:39  */
  assign n11402_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:103:39  */
  assign n11403_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:103:39  */
  assign n11404_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:103:39  */
  assign n11405_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:103:39  */
  assign n11406_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:103:39  */
  assign n11407_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:103:39  */
  assign n11408_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:103:39  */
  assign n11409_o = ci_instr16_i[12];
  assign n11410_o = {n11397_o, n11398_o, n11399_o, n11400_o};
  assign n11411_o = {n11401_o, n11402_o, n11403_o, n11404_o};
  assign n11412_o = {n11405_o, n11406_o, n11407_o, n11408_o};
  assign n11413_o = {n11410_o, n11411_o, n11412_o, n11409_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:105:31  */
  assign n11416_o = ci_instr16_i[3];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:106:31  */
  assign n11418_o = ci_instr16_i[4];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:107:31  */
  assign n11420_o = ci_instr16_i[10];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:108:31  */
  assign n11422_o = ci_instr16_i[11];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:109:31  */
  assign n11424_o = ci_instr16_i[2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:110:31  */
  assign n11426_o = ci_instr16_i[5];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:111:31  */
  assign n11428_o = ci_instr16_i[6];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:112:31  */
  assign n11430_o = ci_instr16_i[12];
  assign n11431_o = n11413_o[12:9];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:22  */
  assign n11432_o = ci_instr16_i[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:26  */
  assign n11433_o = ci_instr16_i[15:13];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:124:87  */
  assign n11436_o = ci_instr16_i[6];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:125:87  */
  assign n11437_o = ci_instr16_i[10];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:126:87  */
  assign n11438_o = ci_instr16_i[11];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:127:87  */
  assign n11439_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:128:87  */
  assign n11440_o = ci_instr16_i[5];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:131:94  */
  assign n11443_o = ci_instr16_i[9:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:131:80  */
  assign n11445_o = {2'b01, n11443_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:132:94  */
  assign n11446_o = ci_instr16_i[4:2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:132:80  */
  assign n11448_o = {2'b01, n11446_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:133:29  */
  assign n11449_o = ci_instr16_i[13];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:133:54  */
  assign n11451_o = n11449_o & 1'b1;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:133:13  */
  assign n11454_o = n11451_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:120:11  */
  assign n11456_o = n11433_o == 3'b010;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:120:22  */
  assign n11458_o = n11433_o == 3'b011;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:120:22  */
  assign n11459_o = n11456_o | n11458_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:141:87  */
  assign n11462_o = ci_instr16_i[6];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:142:87  */
  assign n11463_o = ci_instr16_i[10];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:143:87  */
  assign n11464_o = ci_instr16_i[11];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:144:87  */
  assign n11465_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:145:87  */
  assign n11466_o = ci_instr16_i[5];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:148:94  */
  assign n11469_o = ci_instr16_i[9:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:148:80  */
  assign n11471_o = {2'b01, n11469_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:149:94  */
  assign n11472_o = ci_instr16_i[4:2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:149:80  */
  assign n11474_o = {2'b01, n11472_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:150:29  */
  assign n11475_o = ci_instr16_i[13];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:150:54  */
  assign n11477_o = n11475_o & 1'b1;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:150:13  */
  assign n11480_o = n11477_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:137:11  */
  assign n11482_o = n11433_o == 3'b110;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:137:22  */
  assign n11484_o = n11433_o == 3'b111;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:137:22  */
  assign n11485_o = n11482_o | n11484_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:158:94  */
  assign n11488_o = ci_instr16_i[4:2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:158:80  */
  assign n11490_o = {2'b01, n11488_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:163:87  */
  assign n11497_o = ci_instr16_i[6];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:164:87  */
  assign n11499_o = ci_instr16_i[5];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:165:87  */
  assign n11501_o = ci_instr16_i[11];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:166:87  */
  assign n11503_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:167:87  */
  assign n11505_o = ci_instr16_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:168:87  */
  assign n11507_o = ci_instr16_i[8];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:169:87  */
  assign n11509_o = ci_instr16_i[9];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:170:87  */
  assign n11511_o = ci_instr16_i[10];
  assign n11512_o = n11492_o[11:10];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:172:29  */
  assign n11513_o = ci_instr16_i[12:5];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:172:43  */
  assign n11515_o = n11513_o == 8'b00000000;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:173:29  */
  assign n11516_o = ci_instr16_i[15:13];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:173:70  */
  assign n11518_o = n11516_o == 3'b001;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:172:57  */
  assign n11519_o = n11515_o | n11518_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:174:29  */
  assign n11520_o = ci_instr16_i[15:13];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:174:70  */
  assign n11522_o = n11520_o == 3'b100;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:173:79  */
  assign n11523_o = n11519_o | n11522_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:175:29  */
  assign n11524_o = ci_instr16_i[15:13];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:175:70  */
  assign n11526_o = n11524_o == 3'b101;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:174:79  */
  assign n11527_o = n11523_o | n11526_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:172:13  */
  assign n11530_o = n11527_o ? 1'b1 : 1'b0;
  assign n11531_o = {n11485_o, n11459_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11532_o = n11480_o;
      2'b01: n11532_o = n11454_o;
      default: n11532_o = n11530_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11533_o = 7'b0100011;
      2'b01: n11533_o = 7'b0000011;
      default: n11533_o = 7'b0010011;
    endcase
  assign n11534_o = n11448_o[1:0];
  assign n11535_o = n11490_o[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11536_o = 2'b00;
      2'b01: n11536_o = n11534_o;
      default: n11536_o = n11535_o;
    endcase
  assign n11537_o = n11448_o[2];
  assign n11538_o = n11490_o[2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11539_o = n11462_o;
      2'b01: n11539_o = n11537_o;
      default: n11539_o = n11538_o;
    endcase
  assign n11540_o = n11448_o[3];
  assign n11541_o = n11490_o[3];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11542_o = n11463_o;
      2'b01: n11542_o = n11540_o;
      default: n11542_o = n11541_o;
    endcase
  assign n11543_o = n11448_o[4];
  assign n11544_o = n11490_o[4];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11545_o = n11464_o;
      2'b01: n11545_o = n11543_o;
      default: n11545_o = n11544_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11546_o = 3'b010;
      2'b01: n11546_o = 3'b010;
      default: n11546_o = 3'b000;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11547_o = n11471_o;
      2'b01: n11547_o = n11445_o;
      default: n11547_o = 5'b00010;
    endcase
  assign n11548_o = n11435_o[0];
  assign n11549_o = n11474_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11550_o = n11549_o;
      2'b01: n11550_o = n11548_o;
      default: n11550_o = 1'b0;
    endcase
  assign n11551_o = n11435_o[1];
  assign n11552_o = n11474_o[1];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11553_o = n11552_o;
      2'b01: n11553_o = n11551_o;
      default: n11553_o = 1'b0;
    endcase
  assign n11554_o = n11474_o[2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11555_o = n11554_o;
      2'b01: n11555_o = n11436_o;
      default: n11555_o = n11497_o;
    endcase
  assign n11556_o = n11474_o[3];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11557_o = n11556_o;
      2'b01: n11557_o = n11437_o;
      default: n11557_o = n11499_o;
    endcase
  assign n11558_o = n11474_o[4];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11559_o = n11558_o;
      2'b01: n11559_o = n11438_o;
      default: n11559_o = n11501_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11560_o = n11465_o;
      2'b01: n11560_o = n11439_o;
      default: n11560_o = n11503_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11561_o = n11466_o;
      2'b01: n11561_o = n11440_o;
      default: n11561_o = n11505_o;
    endcase
  assign n11562_o = n11441_o[0];
  assign n11563_o = n11467_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11564_o = n11563_o;
      2'b01: n11564_o = n11562_o;
      default: n11564_o = n11507_o;
    endcase
  assign n11565_o = n11441_o[1];
  assign n11566_o = n11467_o[1];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11567_o = n11566_o;
      2'b01: n11567_o = n11565_o;
      default: n11567_o = n11509_o;
    endcase
  assign n11568_o = n11441_o[2];
  assign n11569_o = n11467_o[2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11570_o = n11569_o;
      2'b01: n11570_o = n11568_o;
      default: n11570_o = n11511_o;
    endcase
  assign n11571_o = n11441_o[4:3];
  assign n11572_o = n11467_o[4:3];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:9  */
  always @*
    case (n11531_o)
      2'b10: n11573_o = n11572_o;
      2'b01: n11573_o = n11571_o;
      default: n11573_o = n11512_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:117:7  */
  assign n11575_o = n11432_o == 2'b00;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:183:26  */
  assign n11576_o = ci_instr16_i[15:13];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:186:29  */
  assign n11577_o = ci_instr16_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:186:13  */
  assign n11580_o = n11577_o ? 5'b00000 : 5'b00001;
  assign n11582_o = {n11396_o, n11395_o, n11393_o, n11391_o, n11389_o, n11387_o, n11385_o, n11383_o, n11381_o, n11379_o, n11377_o, n11375_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:192:82  */
  assign n11583_o = n11582_o[19:12];
  assign n11584_o = {n11396_o, n11395_o, n11393_o, n11391_o, n11389_o, n11387_o, n11385_o, n11383_o, n11381_o, n11379_o, n11377_o, n11375_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:193:82  */
  assign n11585_o = n11584_o[11];
  assign n11586_o = {n11396_o, n11395_o, n11393_o, n11391_o, n11389_o, n11387_o, n11385_o, n11383_o, n11381_o, n11379_o, n11377_o, n11375_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:194:82  */
  assign n11587_o = n11586_o[10:1];
  assign n11588_o = {n11396_o, n11395_o, n11393_o, n11391_o, n11389_o, n11387_o, n11385_o, n11383_o, n11381_o, n11379_o, n11377_o, n11375_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:195:82  */
  assign n11589_o = n11588_o[20];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:184:11  */
  assign n11591_o = n11576_o == 3'b101;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:184:22  */
  assign n11593_o = n11576_o == 3'b001;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:184:22  */
  assign n11594_o = n11591_o | n11593_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:199:29  */
  assign n11595_o = ci_instr16_i[13];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:199:47  */
  assign n11596_o = ~n11595_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:199:13  */
  assign n11599_o = n11596_o ? 3'b000 : 3'b001;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:205:94  */
  assign n11601_o = ci_instr16_i[9:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:205:80  */
  assign n11603_o = {2'b01, n11601_o};
  assign n11605_o = {n11431_o, n11430_o, n11428_o, n11426_o, n11424_o, n11422_o, n11420_o, n11418_o, n11416_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:207:82  */
  assign n11606_o = n11605_o[11];
  assign n11607_o = {n11431_o, n11430_o, n11428_o, n11426_o, n11424_o, n11422_o, n11420_o, n11418_o, n11416_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:208:82  */
  assign n11608_o = n11607_o[4:1];
  assign n11609_o = {n11431_o, n11430_o, n11428_o, n11426_o, n11424_o, n11422_o, n11420_o, n11418_o, n11416_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:209:82  */
  assign n11610_o = n11609_o[10:5];
  assign n11611_o = {n11431_o, n11430_o, n11428_o, n11426_o, n11424_o, n11422_o, n11420_o, n11418_o, n11416_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:210:82  */
  assign n11612_o = n11611_o[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:197:11  */
  assign n11614_o = n11576_o == 3'b110;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:197:22  */
  assign n11616_o = n11576_o == 3'b111;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:197:22  */
  assign n11617_o = n11614_o | n11616_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:217:87  */
  assign n11619_o = ci_instr16_i[11:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:218:98  */
  assign n11620_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:218:98  */
  assign n11621_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:218:98  */
  assign n11622_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:218:98  */
  assign n11623_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:218:98  */
  assign n11624_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:218:98  */
  assign n11625_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:218:98  */
  assign n11626_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:218:98  */
  assign n11627_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:218:98  */
  assign n11628_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:218:98  */
  assign n11629_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:218:98  */
  assign n11630_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:218:98  */
  assign n11631_o = ci_instr16_i[12];
  assign n11632_o = {n11620_o, n11621_o, n11622_o, n11623_o};
  assign n11633_o = {n11624_o, n11625_o, n11626_o, n11627_o};
  assign n11634_o = {n11628_o, n11629_o, n11630_o, n11631_o};
  assign n11635_o = {n11632_o, n11633_o, n11634_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:219:87  */
  assign n11636_o = ci_instr16_i[2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:220:87  */
  assign n11638_o = ci_instr16_i[3];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:221:87  */
  assign n11640_o = ci_instr16_i[4];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:222:87  */
  assign n11642_o = ci_instr16_i[5];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:223:87  */
  assign n11644_o = ci_instr16_i[6];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:224:87  */
  assign n11646_o = ci_instr16_i[12];
  assign n11647_o = n11635_o[11:6];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:212:11  */
  assign n11649_o = n11576_o == 3'b010;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:228:29  */
  assign n11650_o = ci_instr16_i[11:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:228:66  */
  assign n11652_o = n11650_o == 5'b00010;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:234:100  */
  assign n11656_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:234:100  */
  assign n11657_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:234:100  */
  assign n11658_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:234:100  */
  assign n11659_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:234:100  */
  assign n11660_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:234:100  */
  assign n11661_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:234:100  */
  assign n11662_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:234:100  */
  assign n11663_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:234:100  */
  assign n11664_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:234:100  */
  assign n11665_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:234:100  */
  assign n11666_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:234:100  */
  assign n11667_o = ci_instr16_i[12];
  assign n11668_o = {n11656_o, n11657_o, n11658_o, n11659_o};
  assign n11669_o = {n11660_o, n11661_o, n11662_o, n11663_o};
  assign n11670_o = {n11664_o, n11665_o, n11666_o, n11667_o};
  assign n11671_o = {n11668_o, n11669_o, n11670_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:239:89  */
  assign n11680_o = ci_instr16_i[6];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:240:89  */
  assign n11682_o = ci_instr16_i[2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:241:89  */
  assign n11684_o = ci_instr16_i[5];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:242:89  */
  assign n11686_o = ci_instr16_i[3];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:243:89  */
  assign n11688_o = ci_instr16_i[4];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:244:89  */
  assign n11690_o = ci_instr16_i[12];
  assign n11691_o = n11671_o[11:10];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:247:89  */
  assign n11693_o = ci_instr16_i[11:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11694_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11695_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11696_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11697_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11698_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11699_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11700_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11701_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11702_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11703_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11704_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11705_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11706_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11707_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11708_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11709_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11710_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11711_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11712_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:248:100  */
  assign n11713_o = ci_instr16_i[12];
  assign n11714_o = {n11694_o, n11695_o, n11696_o, n11697_o};
  assign n11715_o = {n11698_o, n11699_o, n11700_o, n11701_o};
  assign n11716_o = {n11702_o, n11703_o, n11704_o, n11705_o};
  assign n11717_o = {n11706_o, n11707_o, n11708_o, n11709_o};
  assign n11718_o = {n11710_o, n11711_o, n11712_o, n11713_o};
  assign n11719_o = {n11714_o, n11715_o, n11716_o, n11717_o};
  assign n11720_o = {n11719_o, n11718_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:249:89  */
  assign n11721_o = ci_instr16_i[2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:250:89  */
  assign n11723_o = ci_instr16_i[3];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:251:89  */
  assign n11725_o = ci_instr16_i[4];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:252:89  */
  assign n11727_o = ci_instr16_i[5];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:253:89  */
  assign n11729_o = ci_instr16_i[6];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:254:89  */
  assign n11731_o = ci_instr16_i[12];
  assign n11732_o = n11720_o[19:6];
  assign n11733_o = {n11732_o, n11731_o, n11729_o, n11727_o, n11725_o, n11723_o, n11721_o, n11693_o, 7'b0110111};
  assign n11734_o = {n11691_o, n11690_o, n11688_o, n11686_o, n11684_o, n11682_o, n11680_o, 1'b0, 1'b0, 1'b0, 1'b0, 5'b00010, 3'b000, 5'b00010, 7'b0010011};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:228:13  */
  assign n11735_o = n11652_o ? n11734_o : n11733_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:256:29  */
  assign n11736_o = ci_instr16_i[6:2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:256:42  */
  assign n11738_o = n11736_o == 5'b00000;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:256:70  */
  assign n11739_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:256:75  */
  assign n11740_o = ~n11739_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:256:53  */
  assign n11741_o = n11738_o & n11740_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:256:13  */
  assign n11744_o = n11741_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:226:11  */
  assign n11746_o = n11576_o == 3'b011;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:264:87  */
  assign n11747_o = ci_instr16_i[11:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:265:87  */
  assign n11748_o = ci_instr16_i[11:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:266:98  */
  assign n11749_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:266:98  */
  assign n11750_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:266:98  */
  assign n11751_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:266:98  */
  assign n11752_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:266:98  */
  assign n11753_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:266:98  */
  assign n11754_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:266:98  */
  assign n11755_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:266:98  */
  assign n11756_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:266:98  */
  assign n11757_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:266:98  */
  assign n11758_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:266:98  */
  assign n11759_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:266:98  */
  assign n11760_o = ci_instr16_i[12];
  assign n11761_o = {n11749_o, n11750_o, n11751_o, n11752_o};
  assign n11762_o = {n11753_o, n11754_o, n11755_o, n11756_o};
  assign n11763_o = {n11757_o, n11758_o, n11759_o, n11760_o};
  assign n11764_o = {n11761_o, n11762_o, n11763_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:267:87  */
  assign n11765_o = ci_instr16_i[2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:268:87  */
  assign n11767_o = ci_instr16_i[3];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:269:87  */
  assign n11769_o = ci_instr16_i[4];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:270:87  */
  assign n11771_o = ci_instr16_i[5];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:271:87  */
  assign n11773_o = ci_instr16_i[6];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:272:87  */
  assign n11775_o = ci_instr16_i[12];
  assign n11776_o = n11764_o[11:6];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:260:11  */
  assign n11778_o = n11576_o == 3'b000;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:276:88  */
  assign n11779_o = ci_instr16_i[9:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:276:74  */
  assign n11781_o = {2'b01, n11779_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:277:88  */
  assign n11782_o = ci_instr16_i[9:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:277:74  */
  assign n11784_o = {2'b01, n11782_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:278:88  */
  assign n11785_o = ci_instr16_i[4:2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:278:74  */
  assign n11787_o = {2'b01, n11785_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:279:30  */
  assign n11788_o = ci_instr16_i[11:10];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:281:33  */
  assign n11789_o = ci_instr16_i[10];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:281:38  */
  assign n11790_o = ~n11789_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:281:17  */
  assign n11793_o = n11790_o ? 7'b0000000 : 7'b0100000;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:288:91  */
  assign n11795_o = ci_instr16_i[2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:289:91  */
  assign n11796_o = ci_instr16_i[3];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:290:91  */
  assign n11797_o = ci_instr16_i[4];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:291:91  */
  assign n11798_o = ci_instr16_i[5];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:292:91  */
  assign n11799_o = ci_instr16_i[6];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:293:33  */
  assign n11800_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:293:17  */
  assign n11803_o = n11800_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:280:15  */
  assign n11805_o = n11788_o == 2'b00;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:280:25  */
  assign n11807_o = n11788_o == 2'b01;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:280:25  */
  assign n11808_o = n11805_o | n11807_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:299:102  */
  assign n11810_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:299:102  */
  assign n11811_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:299:102  */
  assign n11812_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:299:102  */
  assign n11813_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:299:102  */
  assign n11814_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:299:102  */
  assign n11815_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:299:102  */
  assign n11816_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:299:102  */
  assign n11817_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:299:102  */
  assign n11818_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:299:102  */
  assign n11819_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:299:102  */
  assign n11820_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:299:102  */
  assign n11821_o = ci_instr16_i[12];
  assign n11822_o = {n11810_o, n11811_o, n11812_o, n11813_o};
  assign n11823_o = {n11814_o, n11815_o, n11816_o, n11817_o};
  assign n11824_o = {n11818_o, n11819_o, n11820_o, n11821_o};
  assign n11825_o = {n11822_o, n11823_o, n11824_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:300:91  */
  assign n11826_o = ci_instr16_i[2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:301:91  */
  assign n11828_o = ci_instr16_i[3];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:302:91  */
  assign n11830_o = ci_instr16_i[4];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:303:91  */
  assign n11832_o = ci_instr16_i[5];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:304:91  */
  assign n11834_o = ci_instr16_i[6];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:305:91  */
  assign n11836_o = ci_instr16_i[12];
  assign n11837_o = n11825_o[11:6];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:296:15  */
  assign n11839_o = n11788_o == 2'b10;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:308:34  */
  assign n11841_o = ci_instr16_i[6:5];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:309:19  */
  assign n11844_o = n11841_o == 2'b00;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:312:19  */
  assign n11848_o = n11841_o == 2'b01;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:315:19  */
  assign n11852_o = n11841_o == 2'b10;
  assign n11854_o = {n11852_o, n11848_o, n11844_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:308:17  */
  always @*
    case (n11854_o)
      3'b100: n11855_o = 3'b110;
      3'b010: n11855_o = 3'b100;
      3'b001: n11855_o = 3'b000;
      default: n11855_o = 3'b111;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:308:17  */
  always @*
    case (n11854_o)
      3'b100: n11856_o = 7'b0000000;
      3'b010: n11856_o = 7'b0000000;
      3'b001: n11856_o = 7'b0100000;
      default: n11856_o = 7'b0000000;
    endcase
  assign n11857_o = {n11839_o, n11808_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:279:13  */
  always @*
    case (n11857_o)
      2'b10: n11859_o = 1'b0;
      2'b01: n11859_o = n11803_o;
      default: n11859_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:279:13  */
  always @*
    case (n11857_o)
      2'b10: n11860_o = 7'b0010011;
      2'b01: n11860_o = 7'b0010011;
      default: n11860_o = 7'b0110011;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:279:13  */
  always @*
    case (n11857_o)
      2'b10: n11861_o = 3'b111;
      2'b01: n11861_o = 3'b101;
      default: n11861_o = n11855_o;
    endcase
  assign n11862_o = n11787_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:279:13  */
  always @*
    case (n11857_o)
      2'b10: n11863_o = n11826_o;
      2'b01: n11863_o = n11795_o;
      default: n11863_o = n11862_o;
    endcase
  assign n11864_o = n11787_o[1];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:279:13  */
  always @*
    case (n11857_o)
      2'b10: n11865_o = n11828_o;
      2'b01: n11865_o = n11796_o;
      default: n11865_o = n11864_o;
    endcase
  assign n11866_o = n11787_o[2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:279:13  */
  always @*
    case (n11857_o)
      2'b10: n11867_o = n11830_o;
      2'b01: n11867_o = n11797_o;
      default: n11867_o = n11866_o;
    endcase
  assign n11868_o = n11787_o[3];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:279:13  */
  always @*
    case (n11857_o)
      2'b10: n11869_o = n11832_o;
      2'b01: n11869_o = n11798_o;
      default: n11869_o = n11868_o;
    endcase
  assign n11870_o = n11787_o[4];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:279:13  */
  always @*
    case (n11857_o)
      2'b10: n11871_o = n11834_o;
      2'b01: n11871_o = n11799_o;
      default: n11871_o = n11870_o;
    endcase
  assign n11872_o = n11793_o[0];
  assign n11873_o = n11856_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:279:13  */
  always @*
    case (n11857_o)
      2'b10: n11874_o = n11836_o;
      2'b01: n11874_o = n11872_o;
      default: n11874_o = n11873_o;
    endcase
  assign n11875_o = n11793_o[6:1];
  assign n11876_o = n11856_o[6:1];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:279:13  */
  always @*
    case (n11857_o)
      2'b10: n11877_o = n11837_o;
      2'b01: n11877_o = n11875_o;
      default: n11877_o = n11876_o;
    endcase
  assign n11882_o = {n11778_o, n11746_o, n11649_o, n11617_o, n11594_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:183:9  */
  always @*
    case (n11882_o)
      5'b10000: n11884_o = 1'b0;
      5'b01000: n11884_o = n11744_o;
      5'b00100: n11884_o = 1'b0;
      5'b00010: n11884_o = 1'b0;
      5'b00001: n11884_o = 1'b0;
      default: n11884_o = n11859_o;
    endcase
  assign n11885_o = n11735_o[6:0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:183:9  */
  always @*
    case (n11882_o)
      5'b10000: n11886_o = 7'b0010011;
      5'b01000: n11886_o = n11885_o;
      5'b00100: n11886_o = 7'b0010011;
      5'b00010: n11886_o = 7'b1100011;
      5'b00001: n11886_o = 7'b1101111;
      default: n11886_o = n11860_o;
    endcase
  assign n11887_o = n11580_o[0];
  assign n11888_o = n11619_o[0];
  assign n11889_o = n11735_o[7];
  assign n11890_o = n11748_o[0];
  assign n11891_o = n11781_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:183:9  */
  always @*
    case (n11882_o)
      5'b10000: n11892_o = n11890_o;
      5'b01000: n11892_o = n11889_o;
      5'b00100: n11892_o = n11888_o;
      5'b00010: n11892_o = n11606_o;
      5'b00001: n11892_o = n11887_o;
      default: n11892_o = n11891_o;
    endcase
  assign n11893_o = n11580_o[4:1];
  assign n11894_o = n11619_o[4:1];
  assign n11895_o = n11735_o[11:8];
  assign n11896_o = n11748_o[4:1];
  assign n11897_o = n11781_o[4:1];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:183:9  */
  always @*
    case (n11882_o)
      5'b10000: n11898_o = n11896_o;
      5'b01000: n11898_o = n11895_o;
      5'b00100: n11898_o = n11894_o;
      5'b00010: n11898_o = n11608_o;
      5'b00001: n11898_o = n11893_o;
      default: n11898_o = n11897_o;
    endcase
  assign n11899_o = n11583_o[2:0];
  assign n11900_o = n11735_o[14:12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:183:9  */
  always @*
    case (n11882_o)
      5'b10000: n11901_o = 3'b000;
      5'b01000: n11901_o = n11900_o;
      5'b00100: n11901_o = 3'b000;
      5'b00010: n11901_o = n11599_o;
      5'b00001: n11901_o = n11899_o;
      default: n11901_o = n11861_o;
    endcase
  assign n11902_o = n11583_o[7:3];
  assign n11903_o = n11735_o[19:15];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:183:9  */
  always @*
    case (n11882_o)
      5'b10000: n11904_o = n11747_o;
      5'b01000: n11904_o = n11903_o;
      5'b00100: n11904_o = 5'b00000;
      5'b00010: n11904_o = n11603_o;
      5'b00001: n11904_o = n11902_o;
      default: n11904_o = n11784_o;
    endcase
  assign n11905_o = n11604_o[0];
  assign n11906_o = n11735_o[20];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:183:9  */
  always @*
    case (n11882_o)
      5'b10000: n11907_o = n11765_o;
      5'b01000: n11907_o = n11906_o;
      5'b00100: n11907_o = n11636_o;
      5'b00010: n11907_o = n11905_o;
      5'b00001: n11907_o = n11585_o;
      default: n11907_o = n11863_o;
    endcase
  assign n11908_o = n11587_o[0];
  assign n11909_o = n11604_o[1];
  assign n11910_o = n11735_o[21];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:183:9  */
  always @*
    case (n11882_o)
      5'b10000: n11911_o = n11767_o;
      5'b01000: n11911_o = n11910_o;
      5'b00100: n11911_o = n11638_o;
      5'b00010: n11911_o = n11909_o;
      5'b00001: n11911_o = n11908_o;
      default: n11911_o = n11865_o;
    endcase
  assign n11912_o = n11587_o[1];
  assign n11913_o = n11604_o[2];
  assign n11914_o = n11735_o[22];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:183:9  */
  always @*
    case (n11882_o)
      5'b10000: n11915_o = n11769_o;
      5'b01000: n11915_o = n11914_o;
      5'b00100: n11915_o = n11640_o;
      5'b00010: n11915_o = n11913_o;
      5'b00001: n11915_o = n11912_o;
      default: n11915_o = n11867_o;
    endcase
  assign n11916_o = n11587_o[2];
  assign n11917_o = n11604_o[3];
  assign n11918_o = n11735_o[23];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:183:9  */
  always @*
    case (n11882_o)
      5'b10000: n11919_o = n11771_o;
      5'b01000: n11919_o = n11918_o;
      5'b00100: n11919_o = n11642_o;
      5'b00010: n11919_o = n11917_o;
      5'b00001: n11919_o = n11916_o;
      default: n11919_o = n11869_o;
    endcase
  assign n11920_o = n11587_o[3];
  assign n11921_o = n11604_o[4];
  assign n11922_o = n11735_o[24];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:183:9  */
  always @*
    case (n11882_o)
      5'b10000: n11923_o = n11773_o;
      5'b01000: n11923_o = n11922_o;
      5'b00100: n11923_o = n11644_o;
      5'b00010: n11923_o = n11921_o;
      5'b00001: n11923_o = n11920_o;
      default: n11923_o = n11871_o;
    endcase
  assign n11924_o = n11587_o[4];
  assign n11925_o = n11610_o[0];
  assign n11926_o = n11735_o[25];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:183:9  */
  always @*
    case (n11882_o)
      5'b10000: n11927_o = n11775_o;
      5'b01000: n11927_o = n11926_o;
      5'b00100: n11927_o = n11646_o;
      5'b00010: n11927_o = n11925_o;
      5'b00001: n11927_o = n11924_o;
      default: n11927_o = n11874_o;
    endcase
  assign n11928_o = n11587_o[9:5];
  assign n11929_o = n11610_o[5:1];
  assign n11930_o = n11647_o[4:0];
  assign n11931_o = n11735_o[30:26];
  assign n11932_o = n11776_o[4:0];
  assign n11933_o = n11877_o[4:0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:183:9  */
  always @*
    case (n11882_o)
      5'b10000: n11934_o = n11932_o;
      5'b01000: n11934_o = n11931_o;
      5'b00100: n11934_o = n11930_o;
      5'b00010: n11934_o = n11929_o;
      5'b00001: n11934_o = n11928_o;
      default: n11934_o = n11933_o;
    endcase
  assign n11935_o = n11647_o[5];
  assign n11936_o = n11735_o[31];
  assign n11937_o = n11776_o[5];
  assign n11938_o = n11877_o[5];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:183:9  */
  always @*
    case (n11882_o)
      5'b10000: n11939_o = n11937_o;
      5'b01000: n11939_o = n11936_o;
      5'b00100: n11939_o = n11935_o;
      5'b00010: n11939_o = n11612_o;
      5'b00001: n11939_o = n11589_o;
      default: n11939_o = n11938_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:181:7  */
  assign n11941_o = n11432_o == 2'b01;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:26  */
  assign n11942_o = ci_instr16_i[15:13];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:332:87  */
  assign n11943_o = ci_instr16_i[11:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:333:87  */
  assign n11944_o = ci_instr16_i[11:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:336:87  */
  assign n11947_o = ci_instr16_i[2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:337:87  */
  assign n11948_o = ci_instr16_i[3];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:338:87  */
  assign n11949_o = ci_instr16_i[4];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:339:87  */
  assign n11950_o = ci_instr16_i[5];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:340:87  */
  assign n11951_o = ci_instr16_i[6];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:341:29  */
  assign n11952_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:341:13  */
  assign n11955_o = n11952_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:329:11  */
  assign n11957_o = n11942_o == 3'b000;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:349:87  */
  assign n11959_o = ci_instr16_i[4];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:350:87  */
  assign n11960_o = ci_instr16_i[5];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:351:87  */
  assign n11961_o = ci_instr16_i[6];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:352:87  */
  assign n11962_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:353:87  */
  assign n11963_o = ci_instr16_i[2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:354:87  */
  assign n11964_o = ci_instr16_i[3];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:358:87  */
  assign n11967_o = ci_instr16_i[11:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:359:29  */
  assign n11968_o = ci_instr16_i[13];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:359:54  */
  assign n11970_o = n11968_o & 1'b1;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:359:13  */
  assign n11973_o = n11970_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:345:11  */
  assign n11975_o = n11942_o == 3'b010;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:345:22  */
  assign n11977_o = n11942_o == 3'b011;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:345:22  */
  assign n11978_o = n11975_o | n11977_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:367:87  */
  assign n11980_o = ci_instr16_i[9];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:368:87  */
  assign n11981_o = ci_instr16_i[10];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:369:87  */
  assign n11982_o = ci_instr16_i[11];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:370:87  */
  assign n11983_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:371:87  */
  assign n11984_o = ci_instr16_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:372:87  */
  assign n11985_o = ci_instr16_i[8];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:376:87  */
  assign n11988_o = ci_instr16_i[6:2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:377:29  */
  assign n11989_o = ci_instr16_i[13];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:377:54  */
  assign n11991_o = n11989_o & 1'b1;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:377:13  */
  assign n11994_o = n11991_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:363:11  */
  assign n11996_o = n11942_o == 3'b110;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:363:22  */
  assign n11998_o = n11942_o == 3'b111;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:363:22  */
  assign n11999_o = n11996_o | n11998_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:383:29  */
  assign n12000_o = ci_instr16_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:383:34  */
  assign n12001_o = ~n12000_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:384:31  */
  assign n12002_o = ci_instr16_i[6:2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:384:44  */
  assign n12004_o = n12002_o == 5'b00000;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:386:91  */
  assign n12006_o = ci_instr16_i[11:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:391:91  */
  assign n12009_o = ci_instr16_i[11:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:393:91  */
  assign n12011_o = ci_instr16_i[6:2];
  assign n12012_o = {n12011_o, 5'b00000, 3'b000, n12009_o, 7'b0110011};
  assign n12013_o = {5'b00000, 7'b1100111};
  assign n12014_o = n12012_o[11:0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:384:15  */
  assign n12015_o = n12004_o ? n12013_o : n12014_o;
  assign n12016_o = n12012_o[14:12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:384:15  */
  assign n12018_o = n12004_o ? 3'b000 : n12016_o;
  assign n12019_o = n12012_o[19:15];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:384:15  */
  assign n12020_o = n12004_o ? n12006_o : n12019_o;
  assign n12021_o = n12012_o[24:20];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:384:15  */
  assign n12023_o = n12004_o ? 5'b00000 : n12021_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:396:31  */
  assign n12024_o = ci_instr16_i[6:2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:396:44  */
  assign n12026_o = n12024_o == 5'b00000;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:397:33  */
  assign n12027_o = ci_instr16_i[11:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:397:47  */
  assign n12029_o = n12027_o == 5'b00000;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:402:93  */
  assign n12032_o = ci_instr16_i[11:7];
  assign n12034_o = {5'b00001, 7'b1100111};
  assign n12035_o = n12034_o[6:0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:397:17  */
  assign n12036_o = n12029_o ? 7'b1110011 : n12035_o;
  assign n12037_o = n12034_o[11:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:397:17  */
  assign n12039_o = n12029_o ? 5'b00000 : n12037_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:397:17  */
  assign n12041_o = n12029_o ? 5'b00000 : n12032_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:397:17  */
  assign n12043_o = n12029_o ? 12'b000000000001 : 12'b000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:408:91  */
  assign n12045_o = ci_instr16_i[11:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:409:91  */
  assign n12046_o = ci_instr16_i[11:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:410:91  */
  assign n12047_o = ci_instr16_i[6:2];
  assign n12048_o = {n12047_o, n12046_o, 3'b000, n12045_o, 7'b0110011};
  assign n12049_o = {n12039_o, n12036_o};
  assign n12050_o = {n12043_o, n12041_o};
  assign n12051_o = n12048_o[11:0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:396:15  */
  assign n12052_o = n12026_o ? n12049_o : n12051_o;
  assign n12053_o = n12048_o[14:12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:396:15  */
  assign n12055_o = n12026_o ? 3'b000 : n12053_o;
  assign n12056_o = n12048_o[24:15];
  assign n12057_o = n12050_o[9:0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:396:15  */
  assign n12058_o = n12026_o ? n12057_o : n12056_o;
  assign n12059_o = n12050_o[16:10];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:396:15  */
  assign n12061_o = n12026_o ? n12059_o : 7'b0000000;
  assign n12062_o = {n12061_o, n12058_o, n12055_o, n12052_o};
  assign n12063_o = {n12023_o, n12020_o, n12018_o, n12015_o};
  assign n12064_o = n12062_o[24:0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:383:13  */
  assign n12065_o = n12001_o ? n12063_o : n12064_o;
  assign n12066_o = n12062_o[31:25];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:383:13  */
  assign n12068_o = n12001_o ? 7'b0000000 : n12066_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:414:29  */
  assign n12069_o = ci_instr16_i[15:13];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:414:70  */
  assign n12071_o = n12069_o == 3'b001;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:415:29  */
  assign n12072_o = ci_instr16_i[15:13];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:415:70  */
  assign n12074_o = n12072_o == 3'b101;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:414:79  */
  assign n12075_o = n12071_o | n12074_o;
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:414:13  */
  assign n12078_o = n12075_o ? 1'b1 : 1'b0;
  assign n12079_o = {n11999_o, n11978_o, n11957_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:9  */
  always @*
    case (n12079_o)
      3'b100: n12080_o = n11994_o;
      3'b010: n12080_o = n11973_o;
      3'b001: n12080_o = n11955_o;
      default: n12080_o = n12078_o;
    endcase
  assign n12081_o = n12065_o[6:0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:9  */
  always @*
    case (n12079_o)
      3'b100: n12082_o = 7'b0100011;
      3'b010: n12082_o = 7'b0000011;
      3'b001: n12082_o = 7'b0010011;
      default: n12082_o = n12081_o;
    endcase
  assign n12083_o = n11944_o[1:0];
  assign n12084_o = n11967_o[1:0];
  assign n12085_o = n12065_o[8:7];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:9  */
  always @*
    case (n12079_o)
      3'b100: n12086_o = 2'b00;
      3'b010: n12086_o = n12084_o;
      3'b001: n12086_o = n12083_o;
      default: n12086_o = n12085_o;
    endcase
  assign n12087_o = n11944_o[2];
  assign n12088_o = n11967_o[2];
  assign n12089_o = n12065_o[9];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:9  */
  always @*
    case (n12079_o)
      3'b100: n12090_o = n11980_o;
      3'b010: n12090_o = n12088_o;
      3'b001: n12090_o = n12087_o;
      default: n12090_o = n12089_o;
    endcase
  assign n12091_o = n11944_o[3];
  assign n12092_o = n11967_o[3];
  assign n12093_o = n12065_o[10];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:9  */
  always @*
    case (n12079_o)
      3'b100: n12094_o = n11981_o;
      3'b010: n12094_o = n12092_o;
      3'b001: n12094_o = n12091_o;
      default: n12094_o = n12093_o;
    endcase
  assign n12095_o = n11944_o[4];
  assign n12096_o = n11967_o[4];
  assign n12097_o = n12065_o[11];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:9  */
  always @*
    case (n12079_o)
      3'b100: n12098_o = n11982_o;
      3'b010: n12098_o = n12096_o;
      3'b001: n12098_o = n12095_o;
      default: n12098_o = n12097_o;
    endcase
  assign n12099_o = n12065_o[14:12];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:9  */
  always @*
    case (n12079_o)
      3'b100: n12100_o = 3'b010;
      3'b010: n12100_o = 3'b010;
      3'b001: n12100_o = 3'b001;
      default: n12100_o = n12099_o;
    endcase
  assign n12101_o = n12065_o[19:15];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:9  */
  always @*
    case (n12079_o)
      3'b100: n12102_o = 5'b00010;
      3'b010: n12102_o = 5'b00010;
      3'b001: n12102_o = n11943_o;
      default: n12102_o = n12101_o;
    endcase
  assign n12103_o = n11958_o[0];
  assign n12104_o = n11988_o[0];
  assign n12105_o = n12065_o[20];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:9  */
  always @*
    case (n12079_o)
      3'b100: n12106_o = n12104_o;
      3'b010: n12106_o = n12103_o;
      3'b001: n12106_o = n11947_o;
      default: n12106_o = n12105_o;
    endcase
  assign n12107_o = n11958_o[1];
  assign n12108_o = n11988_o[1];
  assign n12109_o = n12065_o[21];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:9  */
  always @*
    case (n12079_o)
      3'b100: n12110_o = n12108_o;
      3'b010: n12110_o = n12107_o;
      3'b001: n12110_o = n11948_o;
      default: n12110_o = n12109_o;
    endcase
  assign n12111_o = n11988_o[2];
  assign n12112_o = n12065_o[22];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:9  */
  always @*
    case (n12079_o)
      3'b100: n12113_o = n12111_o;
      3'b010: n12113_o = n11959_o;
      3'b001: n12113_o = n11949_o;
      default: n12113_o = n12112_o;
    endcase
  assign n12114_o = n11988_o[3];
  assign n12115_o = n12065_o[23];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:9  */
  always @*
    case (n12079_o)
      3'b100: n12116_o = n12114_o;
      3'b010: n12116_o = n11960_o;
      3'b001: n12116_o = n11950_o;
      default: n12116_o = n12115_o;
    endcase
  assign n12117_o = n11988_o[4];
  assign n12118_o = n12065_o[24];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:9  */
  always @*
    case (n12079_o)
      3'b100: n12119_o = n12117_o;
      3'b010: n12119_o = n11961_o;
      3'b001: n12119_o = n11951_o;
      default: n12119_o = n12118_o;
    endcase
  assign n12120_o = n11946_o[0];
  assign n12121_o = n12068_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:9  */
  always @*
    case (n12079_o)
      3'b100: n12122_o = n11983_o;
      3'b010: n12122_o = n11962_o;
      3'b001: n12122_o = n12120_o;
      default: n12122_o = n12121_o;
    endcase
  assign n12123_o = n11946_o[1];
  assign n12124_o = n12068_o[1];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:9  */
  always @*
    case (n12079_o)
      3'b100: n12125_o = n11984_o;
      3'b010: n12125_o = n11963_o;
      3'b001: n12125_o = n12123_o;
      default: n12125_o = n12124_o;
    endcase
  assign n12126_o = n11946_o[2];
  assign n12127_o = n12068_o[2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:9  */
  always @*
    case (n12079_o)
      3'b100: n12128_o = n11985_o;
      3'b010: n12128_o = n11964_o;
      3'b001: n12128_o = n12126_o;
      default: n12128_o = n12127_o;
    endcase
  assign n12129_o = n11946_o[6:3];
  assign n12130_o = n12068_o[6:3];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:327:9  */
  always @*
    case (n12079_o)
      3'b100: n12131_o = 4'b0000;
      3'b010: n12131_o = 4'b0000;
      3'b001: n12131_o = n12129_o;
      default: n12131_o = n12130_o;
    endcase
  assign n12132_o = {n11941_o, n11575_o};
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12133_o = n11884_o;
      2'b01: n12133_o = n11532_o;
      default: n12133_o = n12080_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12135_o = n11886_o;
      2'b01: n12135_o = n11533_o;
      default: n12135_o = n12082_o;
    endcase
  assign n12136_o = n11536_o[0];
  assign n12137_o = n12086_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12138_o = n11892_o;
      2'b01: n12138_o = n12136_o;
      default: n12138_o = n12137_o;
    endcase
  assign n12139_o = n11536_o[1];
  assign n12140_o = n11898_o[0];
  assign n12141_o = n12086_o[1];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12142_o = n12140_o;
      2'b01: n12142_o = n12139_o;
      default: n12142_o = n12141_o;
    endcase
  assign n12143_o = n11898_o[1];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12144_o = n12143_o;
      2'b01: n12144_o = n11539_o;
      default: n12144_o = n12090_o;
    endcase
  assign n12145_o = n11898_o[2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12146_o = n12145_o;
      2'b01: n12146_o = n11542_o;
      default: n12146_o = n12094_o;
    endcase
  assign n12147_o = n11898_o[3];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12148_o = n12147_o;
      2'b01: n12148_o = n11545_o;
      default: n12148_o = n12098_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12149_o = n11901_o;
      2'b01: n12149_o = n11546_o;
      default: n12149_o = n12100_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12150_o = n11904_o;
      2'b01: n12150_o = n11547_o;
      default: n12150_o = n12102_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12151_o = n11907_o;
      2'b01: n12151_o = n11550_o;
      default: n12151_o = n12106_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12152_o = n11911_o;
      2'b01: n12152_o = n11553_o;
      default: n12152_o = n12110_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12153_o = n11915_o;
      2'b01: n12153_o = n11555_o;
      default: n12153_o = n12113_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12154_o = n11919_o;
      2'b01: n12154_o = n11557_o;
      default: n12154_o = n12116_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12155_o = n11923_o;
      2'b01: n12155_o = n11559_o;
      default: n12155_o = n12119_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12156_o = n11927_o;
      2'b01: n12156_o = n11560_o;
      default: n12156_o = n12122_o;
    endcase
  assign n12157_o = n11934_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12158_o = n12157_o;
      2'b01: n12158_o = n11561_o;
      default: n12158_o = n12125_o;
    endcase
  assign n12159_o = n11934_o[1];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12160_o = n12159_o;
      2'b01: n12160_o = n11564_o;
      default: n12160_o = n12128_o;
    endcase
  assign n12161_o = n11934_o[2];
  assign n12162_o = n12131_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12163_o = n12161_o;
      2'b01: n12163_o = n11567_o;
      default: n12163_o = n12162_o;
    endcase
  assign n12164_o = n11934_o[3];
  assign n12165_o = n12131_o[1];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12166_o = n12164_o;
      2'b01: n12166_o = n11570_o;
      default: n12166_o = n12165_o;
    endcase
  assign n12167_o = n11573_o[0];
  assign n12168_o = n11934_o[4];
  assign n12169_o = n12131_o[2];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12170_o = n12168_o;
      2'b01: n12170_o = n12167_o;
      default: n12170_o = n12169_o;
    endcase
  assign n12171_o = n11573_o[1];
  assign n12172_o = n12131_o[3];
  /* ../neorv32/rtl/core/neorv32_cpu_decompressor.vhd:115:5  */
  always @*
    case (n12132_o)
      2'b10: n12173_o = n11939_o;
      2'b01: n12173_o = n12171_o;
      default: n12173_o = n12172_o;
    endcase
  assign n12197_o = {n12173_o, n12170_o, n12166_o, n12163_o, n12160_o, n12158_o, n12156_o, n12155_o, n12154_o, n12153_o, n12152_o, n12151_o, n12150_o, n12149_o, n12148_o, n12146_o, n12144_o, n12142_o, n12138_o, n12135_o};
endmodule

module neorv32_fifo_2_18_1489f923c4dca729178b3e3233458550d8dddf29
  (input  clk_i,
   input  rstn_i,
   input  clear_i,
   input  [17:0] wdata_i,
   input  we_i,
   input  re_i,
   output half_o,
   output free_o,
   output [17:0] rdata_o,
   output avail_o);
  wire [65:0] fifo;
  wire [1:0] level_diff;
  wire n11231_o;
  wire n11232_o;
  wire n11233_o;
  wire n11235_o;
  wire n11236_o;
  wire n11237_o;
  wire n11239_o;
  wire n11244_o;
  wire [1:0] n11245_o;
  wire [1:0] n11247_o;
  wire [1:0] n11248_o;
  wire [1:0] n11249_o;
  wire [1:0] n11250_o;
  wire n11252_o;
  wire [1:0] n11253_o;
  wire [1:0] n11255_o;
  wire [1:0] n11256_o;
  wire [1:0] n11257_o;
  wire [1:0] n11258_o;
  wire [3:0] n11259_o;
  wire [3:0] n11262_o;
  wire n11266_o;
  wire n11267_o;
  wire n11268_o;
  wire n11269_o;
  wire n11272_o;
  wire n11273_o;
  wire n11274_o;
  wire n11275_o;
  wire n11276_o;
  wire n11277_o;
  wire n11280_o;
  wire n11281_o;
  wire n11282_o;
  wire n11283_o;
  wire n11284_o;
  wire n11285_o;
  wire [1:0] n11287_o;
  wire [1:0] n11288_o;
  wire [1:0] n11289_o;
  wire n11290_o;
  wire n11291_o;
  wire n11292_o;
  wire n11293_o;
  wire n11294_o;
  wire n11295_o;
  wire n11296_o;
  wire n11297_o;
  wire n11298_o;
  wire n11299_o;
  wire n11302_o;
  wire n11303_o;
  wire n11306_o;
  wire [35:0] n11308_o;
  wire n11317_o;
  wire n11320_o;
  wire [35:0] n11324_o;
  wire [35:0] n11325_o;
  reg [35:0] n11326_q;
  reg [3:0] n11327_q;
  wire [65:0] n11328_o;
  wire n11329_o;
  wire n11330_o;
  wire [17:0] n11331_o;
  wire [17:0] n11332_o;
  wire [17:0] n11333_o;
  wire [17:0] n11334_o;
  wire [35:0] n11335_o;
  wire [17:0] n11336_o;
  wire [17:0] n11337_o;
  wire [17:0] n11338_o;
  assign half_o = n11299_o;
  assign free_o = n11297_o;
  assign rdata_o = n11338_o;
  assign avail_o = n11298_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:84:10  */
  assign fifo = n11328_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:87:10  */
  assign level_diff = n11289_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:99:19  */
  assign n11231_o = 1'b1 ? re_i : n11233_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:99:64  */
  assign n11232_o = fifo[65];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:99:55  */
  assign n11233_o = re_i & n11232_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:100:19  */
  assign n11235_o = 1'b1 ? we_i : n11237_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:100:64  */
  assign n11236_o = fifo[64];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:100:55  */
  assign n11237_o = we_i & n11236_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:107:16  */
  assign n11239_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:114:19  */
  assign n11244_o = fifo[0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:115:55  */
  assign n11245_o = fifo[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:115:62  */
  assign n11247_o = n11245_o + 2'b01;
  assign n11248_o = fifo[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:114:7  */
  assign n11249_o = n11244_o ? n11247_o : n11248_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:112:7  */
  assign n11250_o = clear_i ? 2'b00 : n11249_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:120:19  */
  assign n11252_o = fifo[1];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:121:55  */
  assign n11253_o = fifo[5:4];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:121:62  */
  assign n11255_o = n11253_o + 2'b01;
  assign n11256_o = fifo[5:4];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:120:7  */
  assign n11257_o = n11252_o ? n11255_o : n11256_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:118:7  */
  assign n11258_o = clear_i ? 2'b00 : n11257_o;
  assign n11259_o = {n11258_o, n11250_o};
  assign n11262_o = {2'b00, 2'b00};
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:131:39  */
  assign n11266_o = fifo[4];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:131:80  */
  assign n11267_o = fifo[2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:131:68  */
  assign n11268_o = n11266_o == n11267_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:131:23  */
  assign n11269_o = n11268_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:132:39  */
  assign n11272_o = fifo[5];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:132:70  */
  assign n11273_o = fifo[3];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:132:57  */
  assign n11274_o = n11272_o != n11273_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:132:99  */
  assign n11275_o = fifo[60];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:132:89  */
  assign n11276_o = n11274_o & n11275_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:132:23  */
  assign n11277_o = n11276_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:133:39  */
  assign n11280_o = fifo[5];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:133:70  */
  assign n11281_o = fifo[3];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:133:58  */
  assign n11282_o = n11280_o == n11281_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:133:99  */
  assign n11283_o = fifo[60];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:133:89  */
  assign n11284_o = n11282_o & n11283_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:133:23  */
  assign n11285_o = n11284_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:134:51  */
  assign n11287_o = fifo[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:134:74  */
  assign n11288_o = fifo[5:4];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:134:58  */
  assign n11289_o = n11287_o - n11288_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:135:29  */
  assign n11290_o = level_diff[0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:135:57  */
  assign n11291_o = fifo[62];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:135:49  */
  assign n11292_o = n11290_o | n11291_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:146:26  */
  assign n11293_o = fifo[62];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:146:17  */
  assign n11294_o = ~n11293_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:147:26  */
  assign n11295_o = fifo[61];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:147:17  */
  assign n11296_o = ~n11295_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:154:21  */
  assign n11297_o = fifo[64];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:155:21  */
  assign n11298_o = fifo[65];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:156:21  */
  assign n11299_o = fifo[63];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:183:18  */
  assign n11302_o = fifo[0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:51  */
  assign n11303_o = fifo[2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:21  */
  assign n11306_o = 1'b1 - n11303_o;
  assign n11308_o = fifo[41:6];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:214:60  */
  assign n11317_o = fifo[4];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:214:30  */
  assign n11320_o = 1'b1 - n11317_o;
  assign n11324_o = fifo[41:6];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:182:7  */
  assign n11325_o = n11302_o ? n11335_o : n11324_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:182:7  */
  always @(posedge clk_i)
    n11326_q <= n11325_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:110:5  */
  always @(posedge clk_i or posedge n11239_o)
    if (n11239_o)
      n11327_q <= n11262_o;
    else
      n11327_q <= n11259_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:107:5  */
  assign n11328_o = {n11296_o, n11294_o, n11292_o, n11277_o, n11285_o, n11269_o, 18'b000000000000000000, n11326_q, n11327_q, n11231_o, n11235_o};
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n11329_o = n11306_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n11330_o = ~n11329_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:58:5  */
  assign n11331_o = n11308_o[17:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n11332_o = n11330_o ? wdata_i : n11331_o;
  assign n11333_o = n11308_o[35:18];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n11334_o = n11329_o ? wdata_i : n11333_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:209:5  */
  assign n11335_o = {n11334_o, n11332_o};
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:21  */
  assign n11336_o = fifo[23:6];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n11337_o = fifo[41:24];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:214:29  */
  assign n11338_o = n11320_o ? n11337_o : n11336_o;
endmodule

module neorv32_fifo_256_8_9159cb8bcee7fcb95582f140960cdae72788d326
  (input  clk_i,
   input  rstn_i,
   input  clear_i,
   input  [7:0] wdata_i,
   input  we_i,
   input  re_i,
   output half_o,
   output free_o,
   output [7:0] rdata_o,
   output avail_o);
  wire [2081:0] fifo;
  wire [8:0] level_diff;
  wire n9645_o;
  wire n9646_o;
  wire n9647_o;
  wire n9649_o;
  wire n9650_o;
  wire n9651_o;
  wire n9653_o;
  wire n9658_o;
  wire [8:0] n9659_o;
  wire [8:0] n9661_o;
  wire [8:0] n9662_o;
  wire [8:0] n9663_o;
  wire [8:0] n9664_o;
  wire n9666_o;
  wire [8:0] n9667_o;
  wire [8:0] n9669_o;
  wire [8:0] n9670_o;
  wire [8:0] n9671_o;
  wire [8:0] n9672_o;
  wire [17:0] n9673_o;
  wire [17:0] n9676_o;
  wire [7:0] n9680_o;
  wire [7:0] n9681_o;
  wire n9682_o;
  wire n9683_o;
  wire n9686_o;
  wire n9687_o;
  wire n9688_o;
  wire n9689_o;
  wire n9690_o;
  wire n9691_o;
  wire n9694_o;
  wire n9695_o;
  wire n9696_o;
  wire n9697_o;
  wire n9698_o;
  wire n9699_o;
  wire [8:0] n9701_o;
  wire [8:0] n9702_o;
  wire [8:0] n9703_o;
  wire n9704_o;
  wire n9705_o;
  wire n9706_o;
  wire n9707_o;
  wire n9708_o;
  wire n9709_o;
  wire n9710_o;
  wire n9712_o;
  wire n9714_o;
  wire n9715_o;
  wire n9716_o;
  wire n9729_o;
  wire [7:0] n9730_o;
  wire [7:0] n9733_o;
  wire [2047:0] n9735_o;
  wire [7:0] n9745_o;
  wire [7:0] n9748_o;
  wire [2047:0] n9753_o;
  wire [2047:0] n9754_o;
  reg [2047:0] n9755_q;
  reg [17:0] n9756_q;
  wire [2081:0] n9757_o;
  reg n9758_q;
  reg n9759_q;
  reg [7:0] n9760_q;
  reg n9761_q;
  wire n9762_o;
  wire n9763_o;
  wire n9764_o;
  wire n9765_o;
  wire n9766_o;
  wire n9767_o;
  wire n9768_o;
  wire n9769_o;
  wire n9770_o;
  wire n9771_o;
  wire n9772_o;
  wire n9773_o;
  wire n9774_o;
  wire n9775_o;
  wire n9776_o;
  wire n9777_o;
  wire n9778_o;
  wire n9779_o;
  wire n9780_o;
  wire n9781_o;
  wire n9782_o;
  wire n9783_o;
  wire n9784_o;
  wire n9785_o;
  wire n9786_o;
  wire n9787_o;
  wire n9788_o;
  wire n9789_o;
  wire n9790_o;
  wire n9791_o;
  wire n9792_o;
  wire n9793_o;
  wire n9794_o;
  wire n9795_o;
  wire n9796_o;
  wire n9797_o;
  wire n9798_o;
  wire n9799_o;
  wire n9800_o;
  wire n9801_o;
  wire n9802_o;
  wire n9803_o;
  wire n9804_o;
  wire n9805_o;
  wire n9806_o;
  wire n9807_o;
  wire n9808_o;
  wire n9809_o;
  wire n9810_o;
  wire n9811_o;
  wire n9812_o;
  wire n9813_o;
  wire n9814_o;
  wire n9815_o;
  wire n9816_o;
  wire n9817_o;
  wire n9818_o;
  wire n9819_o;
  wire n9820_o;
  wire n9821_o;
  wire n9822_o;
  wire n9823_o;
  wire n9824_o;
  wire n9825_o;
  wire n9826_o;
  wire n9827_o;
  wire n9828_o;
  wire n9829_o;
  wire n9830_o;
  wire n9831_o;
  wire n9832_o;
  wire n9833_o;
  wire n9834_o;
  wire n9835_o;
  wire n9836_o;
  wire n9837_o;
  wire n9838_o;
  wire n9839_o;
  wire n9840_o;
  wire n9841_o;
  wire n9842_o;
  wire n9843_o;
  wire n9844_o;
  wire n9845_o;
  wire n9846_o;
  wire n9847_o;
  wire n9848_o;
  wire n9849_o;
  wire n9850_o;
  wire n9851_o;
  wire n9852_o;
  wire n9853_o;
  wire n9854_o;
  wire n9855_o;
  wire n9856_o;
  wire n9857_o;
  wire n9858_o;
  wire n9859_o;
  wire n9860_o;
  wire n9861_o;
  wire n9862_o;
  wire n9863_o;
  wire n9864_o;
  wire n9865_o;
  wire n9866_o;
  wire n9867_o;
  wire n9868_o;
  wire n9869_o;
  wire n9870_o;
  wire n9871_o;
  wire n9872_o;
  wire n9873_o;
  wire n9874_o;
  wire n9875_o;
  wire n9876_o;
  wire n9877_o;
  wire n9878_o;
  wire n9879_o;
  wire n9880_o;
  wire n9881_o;
  wire n9882_o;
  wire n9883_o;
  wire n9884_o;
  wire n9885_o;
  wire n9886_o;
  wire n9887_o;
  wire n9888_o;
  wire n9889_o;
  wire n9890_o;
  wire n9891_o;
  wire n9892_o;
  wire n9893_o;
  wire n9894_o;
  wire n9895_o;
  wire n9896_o;
  wire n9897_o;
  wire n9898_o;
  wire n9899_o;
  wire n9900_o;
  wire n9901_o;
  wire n9902_o;
  wire n9903_o;
  wire n9904_o;
  wire n9905_o;
  wire n9906_o;
  wire n9907_o;
  wire n9908_o;
  wire n9909_o;
  wire n9910_o;
  wire n9911_o;
  wire n9912_o;
  wire n9913_o;
  wire n9914_o;
  wire n9915_o;
  wire n9916_o;
  wire n9917_o;
  wire n9918_o;
  wire n9919_o;
  wire n9920_o;
  wire n9921_o;
  wire n9922_o;
  wire n9923_o;
  wire n9924_o;
  wire n9925_o;
  wire n9926_o;
  wire n9927_o;
  wire n9928_o;
  wire n9929_o;
  wire n9930_o;
  wire n9931_o;
  wire n9932_o;
  wire n9933_o;
  wire n9934_o;
  wire n9935_o;
  wire n9936_o;
  wire n9937_o;
  wire n9938_o;
  wire n9939_o;
  wire n9940_o;
  wire n9941_o;
  wire n9942_o;
  wire n9943_o;
  wire n9944_o;
  wire n9945_o;
  wire n9946_o;
  wire n9947_o;
  wire n9948_o;
  wire n9949_o;
  wire n9950_o;
  wire n9951_o;
  wire n9952_o;
  wire n9953_o;
  wire n9954_o;
  wire n9955_o;
  wire n9956_o;
  wire n9957_o;
  wire n9958_o;
  wire n9959_o;
  wire n9960_o;
  wire n9961_o;
  wire n9962_o;
  wire n9963_o;
  wire n9964_o;
  wire n9965_o;
  wire n9966_o;
  wire n9967_o;
  wire n9968_o;
  wire n9969_o;
  wire n9970_o;
  wire n9971_o;
  wire n9972_o;
  wire n9973_o;
  wire n9974_o;
  wire n9975_o;
  wire n9976_o;
  wire n9977_o;
  wire n9978_o;
  wire n9979_o;
  wire n9980_o;
  wire n9981_o;
  wire n9982_o;
  wire n9983_o;
  wire n9984_o;
  wire n9985_o;
  wire n9986_o;
  wire n9987_o;
  wire n9988_o;
  wire n9989_o;
  wire n9990_o;
  wire n9991_o;
  wire n9992_o;
  wire n9993_o;
  wire n9994_o;
  wire n9995_o;
  wire n9996_o;
  wire n9997_o;
  wire n9998_o;
  wire n9999_o;
  wire n10000_o;
  wire n10001_o;
  wire n10002_o;
  wire n10003_o;
  wire n10004_o;
  wire n10005_o;
  wire n10006_o;
  wire n10007_o;
  wire n10008_o;
  wire n10009_o;
  wire n10010_o;
  wire n10011_o;
  wire n10012_o;
  wire n10013_o;
  wire n10014_o;
  wire n10015_o;
  wire n10016_o;
  wire n10017_o;
  wire n10018_o;
  wire n10019_o;
  wire n10020_o;
  wire n10021_o;
  wire n10022_o;
  wire n10023_o;
  wire n10024_o;
  wire n10025_o;
  wire n10026_o;
  wire n10027_o;
  wire n10028_o;
  wire n10029_o;
  wire n10030_o;
  wire n10031_o;
  wire n10032_o;
  wire n10033_o;
  wire n10034_o;
  wire n10035_o;
  wire n10036_o;
  wire n10037_o;
  wire n10038_o;
  wire n10039_o;
  wire n10040_o;
  wire n10041_o;
  wire n10042_o;
  wire n10043_o;
  wire n10044_o;
  wire n10045_o;
  wire n10046_o;
  wire n10047_o;
  wire n10048_o;
  wire n10049_o;
  wire n10050_o;
  wire n10051_o;
  wire n10052_o;
  wire n10053_o;
  wire n10054_o;
  wire n10055_o;
  wire n10056_o;
  wire n10057_o;
  wire n10058_o;
  wire n10059_o;
  wire n10060_o;
  wire n10061_o;
  wire n10062_o;
  wire n10063_o;
  wire n10064_o;
  wire n10065_o;
  wire n10066_o;
  wire n10067_o;
  wire n10068_o;
  wire n10069_o;
  wire n10070_o;
  wire n10071_o;
  wire n10072_o;
  wire n10073_o;
  wire n10074_o;
  wire n10075_o;
  wire n10076_o;
  wire n10077_o;
  wire n10078_o;
  wire n10079_o;
  wire n10080_o;
  wire n10081_o;
  wire n10082_o;
  wire n10083_o;
  wire n10084_o;
  wire n10085_o;
  wire n10086_o;
  wire n10087_o;
  wire n10088_o;
  wire n10089_o;
  wire n10090_o;
  wire n10091_o;
  wire n10092_o;
  wire n10093_o;
  wire n10094_o;
  wire n10095_o;
  wire n10096_o;
  wire n10097_o;
  wire n10098_o;
  wire n10099_o;
  wire n10100_o;
  wire n10101_o;
  wire n10102_o;
  wire n10103_o;
  wire n10104_o;
  wire n10105_o;
  wire n10106_o;
  wire n10107_o;
  wire n10108_o;
  wire n10109_o;
  wire n10110_o;
  wire n10111_o;
  wire n10112_o;
  wire n10113_o;
  wire n10114_o;
  wire n10115_o;
  wire n10116_o;
  wire n10117_o;
  wire n10118_o;
  wire n10119_o;
  wire n10120_o;
  wire n10121_o;
  wire n10122_o;
  wire n10123_o;
  wire n10124_o;
  wire n10125_o;
  wire n10126_o;
  wire n10127_o;
  wire n10128_o;
  wire n10129_o;
  wire n10130_o;
  wire n10131_o;
  wire n10132_o;
  wire n10133_o;
  wire n10134_o;
  wire n10135_o;
  wire n10136_o;
  wire n10137_o;
  wire n10138_o;
  wire n10139_o;
  wire n10140_o;
  wire n10141_o;
  wire n10142_o;
  wire n10143_o;
  wire n10144_o;
  wire n10145_o;
  wire n10146_o;
  wire n10147_o;
  wire n10148_o;
  wire n10149_o;
  wire n10150_o;
  wire n10151_o;
  wire n10152_o;
  wire n10153_o;
  wire n10154_o;
  wire n10155_o;
  wire n10156_o;
  wire n10157_o;
  wire n10158_o;
  wire n10159_o;
  wire n10160_o;
  wire n10161_o;
  wire n10162_o;
  wire n10163_o;
  wire n10164_o;
  wire n10165_o;
  wire n10166_o;
  wire n10167_o;
  wire n10168_o;
  wire n10169_o;
  wire n10170_o;
  wire n10171_o;
  wire n10172_o;
  wire n10173_o;
  wire n10174_o;
  wire n10175_o;
  wire n10176_o;
  wire n10177_o;
  wire n10178_o;
  wire n10179_o;
  wire n10180_o;
  wire n10181_o;
  wire n10182_o;
  wire n10183_o;
  wire n10184_o;
  wire n10185_o;
  wire n10186_o;
  wire n10187_o;
  wire n10188_o;
  wire n10189_o;
  wire n10190_o;
  wire n10191_o;
  wire n10192_o;
  wire n10193_o;
  wire n10194_o;
  wire n10195_o;
  wire n10196_o;
  wire n10197_o;
  wire n10198_o;
  wire n10199_o;
  wire n10200_o;
  wire n10201_o;
  wire n10202_o;
  wire n10203_o;
  wire n10204_o;
  wire n10205_o;
  wire n10206_o;
  wire n10207_o;
  wire n10208_o;
  wire n10209_o;
  wire n10210_o;
  wire n10211_o;
  wire n10212_o;
  wire n10213_o;
  wire n10214_o;
  wire n10215_o;
  wire n10216_o;
  wire n10217_o;
  wire n10218_o;
  wire n10219_o;
  wire n10220_o;
  wire n10221_o;
  wire n10222_o;
  wire n10223_o;
  wire n10224_o;
  wire n10225_o;
  wire n10226_o;
  wire n10227_o;
  wire n10228_o;
  wire n10229_o;
  wire n10230_o;
  wire n10231_o;
  wire n10232_o;
  wire n10233_o;
  wire n10234_o;
  wire n10235_o;
  wire n10236_o;
  wire n10237_o;
  wire n10238_o;
  wire n10239_o;
  wire n10240_o;
  wire n10241_o;
  wire n10242_o;
  wire n10243_o;
  wire n10244_o;
  wire n10245_o;
  wire n10246_o;
  wire n10247_o;
  wire n10248_o;
  wire n10249_o;
  wire n10250_o;
  wire n10251_o;
  wire n10252_o;
  wire n10253_o;
  wire n10254_o;
  wire n10255_o;
  wire n10256_o;
  wire n10257_o;
  wire n10258_o;
  wire n10259_o;
  wire n10260_o;
  wire n10261_o;
  wire n10262_o;
  wire n10263_o;
  wire n10264_o;
  wire n10265_o;
  wire n10266_o;
  wire n10267_o;
  wire n10268_o;
  wire n10269_o;
  wire n10270_o;
  wire n10271_o;
  wire n10272_o;
  wire n10273_o;
  wire n10274_o;
  wire n10275_o;
  wire n10276_o;
  wire n10277_o;
  wire n10278_o;
  wire n10279_o;
  wire n10280_o;
  wire n10281_o;
  wire n10282_o;
  wire n10283_o;
  wire n10284_o;
  wire n10285_o;
  wire [7:0] n10286_o;
  wire [7:0] n10287_o;
  wire [7:0] n10288_o;
  wire [7:0] n10289_o;
  wire [7:0] n10290_o;
  wire [7:0] n10291_o;
  wire [7:0] n10292_o;
  wire [7:0] n10293_o;
  wire [7:0] n10294_o;
  wire [7:0] n10295_o;
  wire [7:0] n10296_o;
  wire [7:0] n10297_o;
  wire [7:0] n10298_o;
  wire [7:0] n10299_o;
  wire [7:0] n10300_o;
  wire [7:0] n10301_o;
  wire [7:0] n10302_o;
  wire [7:0] n10303_o;
  wire [7:0] n10304_o;
  wire [7:0] n10305_o;
  wire [7:0] n10306_o;
  wire [7:0] n10307_o;
  wire [7:0] n10308_o;
  wire [7:0] n10309_o;
  wire [7:0] n10310_o;
  wire [7:0] n10311_o;
  wire [7:0] n10312_o;
  wire [7:0] n10313_o;
  wire [7:0] n10314_o;
  wire [7:0] n10315_o;
  wire [7:0] n10316_o;
  wire [7:0] n10317_o;
  wire [7:0] n10318_o;
  wire [7:0] n10319_o;
  wire [7:0] n10320_o;
  wire [7:0] n10321_o;
  wire [7:0] n10322_o;
  wire [7:0] n10323_o;
  wire [7:0] n10324_o;
  wire [7:0] n10325_o;
  wire [7:0] n10326_o;
  wire [7:0] n10327_o;
  wire [7:0] n10328_o;
  wire [7:0] n10329_o;
  wire [7:0] n10330_o;
  wire [7:0] n10331_o;
  wire [7:0] n10332_o;
  wire [7:0] n10333_o;
  wire [7:0] n10334_o;
  wire [7:0] n10335_o;
  wire [7:0] n10336_o;
  wire [7:0] n10337_o;
  wire [7:0] n10338_o;
  wire [7:0] n10339_o;
  wire [7:0] n10340_o;
  wire [7:0] n10341_o;
  wire [7:0] n10342_o;
  wire [7:0] n10343_o;
  wire [7:0] n10344_o;
  wire [7:0] n10345_o;
  wire [7:0] n10346_o;
  wire [7:0] n10347_o;
  wire [7:0] n10348_o;
  wire [7:0] n10349_o;
  wire [7:0] n10350_o;
  wire [7:0] n10351_o;
  wire [7:0] n10352_o;
  wire [7:0] n10353_o;
  wire [7:0] n10354_o;
  wire [7:0] n10355_o;
  wire [7:0] n10356_o;
  wire [7:0] n10357_o;
  wire [7:0] n10358_o;
  wire [7:0] n10359_o;
  wire [7:0] n10360_o;
  wire [7:0] n10361_o;
  wire [7:0] n10362_o;
  wire [7:0] n10363_o;
  wire [7:0] n10364_o;
  wire [7:0] n10365_o;
  wire [7:0] n10366_o;
  wire [7:0] n10367_o;
  wire [7:0] n10368_o;
  wire [7:0] n10369_o;
  wire [7:0] n10370_o;
  wire [7:0] n10371_o;
  wire [7:0] n10372_o;
  wire [7:0] n10373_o;
  wire [7:0] n10374_o;
  wire [7:0] n10375_o;
  wire [7:0] n10376_o;
  wire [7:0] n10377_o;
  wire [7:0] n10378_o;
  wire [7:0] n10379_o;
  wire [7:0] n10380_o;
  wire [7:0] n10381_o;
  wire [7:0] n10382_o;
  wire [7:0] n10383_o;
  wire [7:0] n10384_o;
  wire [7:0] n10385_o;
  wire [7:0] n10386_o;
  wire [7:0] n10387_o;
  wire [7:0] n10388_o;
  wire [7:0] n10389_o;
  wire [7:0] n10390_o;
  wire [7:0] n10391_o;
  wire [7:0] n10392_o;
  wire [7:0] n10393_o;
  wire [7:0] n10394_o;
  wire [7:0] n10395_o;
  wire [7:0] n10396_o;
  wire [7:0] n10397_o;
  wire [7:0] n10398_o;
  wire [7:0] n10399_o;
  wire [7:0] n10400_o;
  wire [7:0] n10401_o;
  wire [7:0] n10402_o;
  wire [7:0] n10403_o;
  wire [7:0] n10404_o;
  wire [7:0] n10405_o;
  wire [7:0] n10406_o;
  wire [7:0] n10407_o;
  wire [7:0] n10408_o;
  wire [7:0] n10409_o;
  wire [7:0] n10410_o;
  wire [7:0] n10411_o;
  wire [7:0] n10412_o;
  wire [7:0] n10413_o;
  wire [7:0] n10414_o;
  wire [7:0] n10415_o;
  wire [7:0] n10416_o;
  wire [7:0] n10417_o;
  wire [7:0] n10418_o;
  wire [7:0] n10419_o;
  wire [7:0] n10420_o;
  wire [7:0] n10421_o;
  wire [7:0] n10422_o;
  wire [7:0] n10423_o;
  wire [7:0] n10424_o;
  wire [7:0] n10425_o;
  wire [7:0] n10426_o;
  wire [7:0] n10427_o;
  wire [7:0] n10428_o;
  wire [7:0] n10429_o;
  wire [7:0] n10430_o;
  wire [7:0] n10431_o;
  wire [7:0] n10432_o;
  wire [7:0] n10433_o;
  wire [7:0] n10434_o;
  wire [7:0] n10435_o;
  wire [7:0] n10436_o;
  wire [7:0] n10437_o;
  wire [7:0] n10438_o;
  wire [7:0] n10439_o;
  wire [7:0] n10440_o;
  wire [7:0] n10441_o;
  wire [7:0] n10442_o;
  wire [7:0] n10443_o;
  wire [7:0] n10444_o;
  wire [7:0] n10445_o;
  wire [7:0] n10446_o;
  wire [7:0] n10447_o;
  wire [7:0] n10448_o;
  wire [7:0] n10449_o;
  wire [7:0] n10450_o;
  wire [7:0] n10451_o;
  wire [7:0] n10452_o;
  wire [7:0] n10453_o;
  wire [7:0] n10454_o;
  wire [7:0] n10455_o;
  wire [7:0] n10456_o;
  wire [7:0] n10457_o;
  wire [7:0] n10458_o;
  wire [7:0] n10459_o;
  wire [7:0] n10460_o;
  wire [7:0] n10461_o;
  wire [7:0] n10462_o;
  wire [7:0] n10463_o;
  wire [7:0] n10464_o;
  wire [7:0] n10465_o;
  wire [7:0] n10466_o;
  wire [7:0] n10467_o;
  wire [7:0] n10468_o;
  wire [7:0] n10469_o;
  wire [7:0] n10470_o;
  wire [7:0] n10471_o;
  wire [7:0] n10472_o;
  wire [7:0] n10473_o;
  wire [7:0] n10474_o;
  wire [7:0] n10475_o;
  wire [7:0] n10476_o;
  wire [7:0] n10477_o;
  wire [7:0] n10478_o;
  wire [7:0] n10479_o;
  wire [7:0] n10480_o;
  wire [7:0] n10481_o;
  wire [7:0] n10482_o;
  wire [7:0] n10483_o;
  wire [7:0] n10484_o;
  wire [7:0] n10485_o;
  wire [7:0] n10486_o;
  wire [7:0] n10487_o;
  wire [7:0] n10488_o;
  wire [7:0] n10489_o;
  wire [7:0] n10490_o;
  wire [7:0] n10491_o;
  wire [7:0] n10492_o;
  wire [7:0] n10493_o;
  wire [7:0] n10494_o;
  wire [7:0] n10495_o;
  wire [7:0] n10496_o;
  wire [7:0] n10497_o;
  wire [7:0] n10498_o;
  wire [7:0] n10499_o;
  wire [7:0] n10500_o;
  wire [7:0] n10501_o;
  wire [7:0] n10502_o;
  wire [7:0] n10503_o;
  wire [7:0] n10504_o;
  wire [7:0] n10505_o;
  wire [7:0] n10506_o;
  wire [7:0] n10507_o;
  wire [7:0] n10508_o;
  wire [7:0] n10509_o;
  wire [7:0] n10510_o;
  wire [7:0] n10511_o;
  wire [7:0] n10512_o;
  wire [7:0] n10513_o;
  wire [7:0] n10514_o;
  wire [7:0] n10515_o;
  wire [7:0] n10516_o;
  wire [7:0] n10517_o;
  wire [7:0] n10518_o;
  wire [7:0] n10519_o;
  wire [7:0] n10520_o;
  wire [7:0] n10521_o;
  wire [7:0] n10522_o;
  wire [7:0] n10523_o;
  wire [7:0] n10524_o;
  wire [7:0] n10525_o;
  wire [7:0] n10526_o;
  wire [7:0] n10527_o;
  wire [7:0] n10528_o;
  wire [7:0] n10529_o;
  wire [7:0] n10530_o;
  wire [7:0] n10531_o;
  wire [7:0] n10532_o;
  wire [7:0] n10533_o;
  wire [7:0] n10534_o;
  wire [7:0] n10535_o;
  wire [7:0] n10536_o;
  wire [7:0] n10537_o;
  wire [7:0] n10538_o;
  wire [7:0] n10539_o;
  wire [7:0] n10540_o;
  wire [7:0] n10541_o;
  wire [7:0] n10542_o;
  wire [7:0] n10543_o;
  wire [7:0] n10544_o;
  wire [7:0] n10545_o;
  wire [7:0] n10546_o;
  wire [7:0] n10547_o;
  wire [7:0] n10548_o;
  wire [7:0] n10549_o;
  wire [7:0] n10550_o;
  wire [7:0] n10551_o;
  wire [7:0] n10552_o;
  wire [7:0] n10553_o;
  wire [7:0] n10554_o;
  wire [7:0] n10555_o;
  wire [7:0] n10556_o;
  wire [7:0] n10557_o;
  wire [7:0] n10558_o;
  wire [7:0] n10559_o;
  wire [7:0] n10560_o;
  wire [7:0] n10561_o;
  wire [7:0] n10562_o;
  wire [7:0] n10563_o;
  wire [7:0] n10564_o;
  wire [7:0] n10565_o;
  wire [7:0] n10566_o;
  wire [7:0] n10567_o;
  wire [7:0] n10568_o;
  wire [7:0] n10569_o;
  wire [7:0] n10570_o;
  wire [7:0] n10571_o;
  wire [7:0] n10572_o;
  wire [7:0] n10573_o;
  wire [7:0] n10574_o;
  wire [7:0] n10575_o;
  wire [7:0] n10576_o;
  wire [7:0] n10577_o;
  wire [7:0] n10578_o;
  wire [7:0] n10579_o;
  wire [7:0] n10580_o;
  wire [7:0] n10581_o;
  wire [7:0] n10582_o;
  wire [7:0] n10583_o;
  wire [7:0] n10584_o;
  wire [7:0] n10585_o;
  wire [7:0] n10586_o;
  wire [7:0] n10587_o;
  wire [7:0] n10588_o;
  wire [7:0] n10589_o;
  wire [7:0] n10590_o;
  wire [7:0] n10591_o;
  wire [7:0] n10592_o;
  wire [7:0] n10593_o;
  wire [7:0] n10594_o;
  wire [7:0] n10595_o;
  wire [7:0] n10596_o;
  wire [7:0] n10597_o;
  wire [7:0] n10598_o;
  wire [7:0] n10599_o;
  wire [7:0] n10600_o;
  wire [7:0] n10601_o;
  wire [7:0] n10602_o;
  wire [7:0] n10603_o;
  wire [7:0] n10604_o;
  wire [7:0] n10605_o;
  wire [7:0] n10606_o;
  wire [7:0] n10607_o;
  wire [7:0] n10608_o;
  wire [7:0] n10609_o;
  wire [7:0] n10610_o;
  wire [7:0] n10611_o;
  wire [7:0] n10612_o;
  wire [7:0] n10613_o;
  wire [7:0] n10614_o;
  wire [7:0] n10615_o;
  wire [7:0] n10616_o;
  wire [7:0] n10617_o;
  wire [7:0] n10618_o;
  wire [7:0] n10619_o;
  wire [7:0] n10620_o;
  wire [7:0] n10621_o;
  wire [7:0] n10622_o;
  wire [7:0] n10623_o;
  wire [7:0] n10624_o;
  wire [7:0] n10625_o;
  wire [7:0] n10626_o;
  wire [7:0] n10627_o;
  wire [7:0] n10628_o;
  wire [7:0] n10629_o;
  wire [7:0] n10630_o;
  wire [7:0] n10631_o;
  wire [7:0] n10632_o;
  wire [7:0] n10633_o;
  wire [7:0] n10634_o;
  wire [7:0] n10635_o;
  wire [7:0] n10636_o;
  wire [7:0] n10637_o;
  wire [7:0] n10638_o;
  wire [7:0] n10639_o;
  wire [7:0] n10640_o;
  wire [7:0] n10641_o;
  wire [7:0] n10642_o;
  wire [7:0] n10643_o;
  wire [7:0] n10644_o;
  wire [7:0] n10645_o;
  wire [7:0] n10646_o;
  wire [7:0] n10647_o;
  wire [7:0] n10648_o;
  wire [7:0] n10649_o;
  wire [7:0] n10650_o;
  wire [7:0] n10651_o;
  wire [7:0] n10652_o;
  wire [7:0] n10653_o;
  wire [7:0] n10654_o;
  wire [7:0] n10655_o;
  wire [7:0] n10656_o;
  wire [7:0] n10657_o;
  wire [7:0] n10658_o;
  wire [7:0] n10659_o;
  wire [7:0] n10660_o;
  wire [7:0] n10661_o;
  wire [7:0] n10662_o;
  wire [7:0] n10663_o;
  wire [7:0] n10664_o;
  wire [7:0] n10665_o;
  wire [7:0] n10666_o;
  wire [7:0] n10667_o;
  wire [7:0] n10668_o;
  wire [7:0] n10669_o;
  wire [7:0] n10670_o;
  wire [7:0] n10671_o;
  wire [7:0] n10672_o;
  wire [7:0] n10673_o;
  wire [7:0] n10674_o;
  wire [7:0] n10675_o;
  wire [7:0] n10676_o;
  wire [7:0] n10677_o;
  wire [7:0] n10678_o;
  wire [7:0] n10679_o;
  wire [7:0] n10680_o;
  wire [7:0] n10681_o;
  wire [7:0] n10682_o;
  wire [7:0] n10683_o;
  wire [7:0] n10684_o;
  wire [7:0] n10685_o;
  wire [7:0] n10686_o;
  wire [7:0] n10687_o;
  wire [7:0] n10688_o;
  wire [7:0] n10689_o;
  wire [7:0] n10690_o;
  wire [7:0] n10691_o;
  wire [7:0] n10692_o;
  wire [7:0] n10693_o;
  wire [7:0] n10694_o;
  wire [7:0] n10695_o;
  wire [7:0] n10696_o;
  wire [7:0] n10697_o;
  wire [7:0] n10698_o;
  wire [7:0] n10699_o;
  wire [7:0] n10700_o;
  wire [7:0] n10701_o;
  wire [7:0] n10702_o;
  wire [7:0] n10703_o;
  wire [7:0] n10704_o;
  wire [7:0] n10705_o;
  wire [7:0] n10706_o;
  wire [7:0] n10707_o;
  wire [7:0] n10708_o;
  wire [7:0] n10709_o;
  wire [7:0] n10710_o;
  wire [7:0] n10711_o;
  wire [7:0] n10712_o;
  wire [7:0] n10713_o;
  wire [7:0] n10714_o;
  wire [7:0] n10715_o;
  wire [7:0] n10716_o;
  wire [7:0] n10717_o;
  wire [7:0] n10718_o;
  wire [7:0] n10719_o;
  wire [7:0] n10720_o;
  wire [7:0] n10721_o;
  wire [7:0] n10722_o;
  wire [7:0] n10723_o;
  wire [7:0] n10724_o;
  wire [7:0] n10725_o;
  wire [7:0] n10726_o;
  wire [7:0] n10727_o;
  wire [7:0] n10728_o;
  wire [7:0] n10729_o;
  wire [7:0] n10730_o;
  wire [7:0] n10731_o;
  wire [7:0] n10732_o;
  wire [7:0] n10733_o;
  wire [7:0] n10734_o;
  wire [7:0] n10735_o;
  wire [7:0] n10736_o;
  wire [7:0] n10737_o;
  wire [7:0] n10738_o;
  wire [7:0] n10739_o;
  wire [7:0] n10740_o;
  wire [7:0] n10741_o;
  wire [7:0] n10742_o;
  wire [7:0] n10743_o;
  wire [7:0] n10744_o;
  wire [7:0] n10745_o;
  wire [7:0] n10746_o;
  wire [7:0] n10747_o;
  wire [7:0] n10748_o;
  wire [7:0] n10749_o;
  wire [7:0] n10750_o;
  wire [7:0] n10751_o;
  wire [7:0] n10752_o;
  wire [7:0] n10753_o;
  wire [7:0] n10754_o;
  wire [7:0] n10755_o;
  wire [7:0] n10756_o;
  wire [7:0] n10757_o;
  wire [7:0] n10758_o;
  wire [7:0] n10759_o;
  wire [7:0] n10760_o;
  wire [7:0] n10761_o;
  wire [7:0] n10762_o;
  wire [7:0] n10763_o;
  wire [7:0] n10764_o;
  wire [7:0] n10765_o;
  wire [7:0] n10766_o;
  wire [7:0] n10767_o;
  wire [7:0] n10768_o;
  wire [7:0] n10769_o;
  wire [7:0] n10770_o;
  wire [7:0] n10771_o;
  wire [7:0] n10772_o;
  wire [7:0] n10773_o;
  wire [7:0] n10774_o;
  wire [7:0] n10775_o;
  wire [7:0] n10776_o;
  wire [7:0] n10777_o;
  wire [7:0] n10778_o;
  wire [7:0] n10779_o;
  wire [7:0] n10780_o;
  wire [7:0] n10781_o;
  wire [7:0] n10782_o;
  wire [7:0] n10783_o;
  wire [7:0] n10784_o;
  wire [7:0] n10785_o;
  wire [7:0] n10786_o;
  wire [7:0] n10787_o;
  wire [7:0] n10788_o;
  wire [7:0] n10789_o;
  wire [7:0] n10790_o;
  wire [7:0] n10791_o;
  wire [7:0] n10792_o;
  wire [7:0] n10793_o;
  wire [7:0] n10794_o;
  wire [7:0] n10795_o;
  wire [7:0] n10796_o;
  wire [7:0] n10797_o;
  wire [2047:0] n10798_o;
  wire [7:0] n10799_o;
  wire [7:0] n10800_o;
  wire [7:0] n10801_o;
  wire [7:0] n10802_o;
  wire [7:0] n10803_o;
  wire [7:0] n10804_o;
  wire [7:0] n10805_o;
  wire [7:0] n10806_o;
  wire [7:0] n10807_o;
  wire [7:0] n10808_o;
  wire [7:0] n10809_o;
  wire [7:0] n10810_o;
  wire [7:0] n10811_o;
  wire [7:0] n10812_o;
  wire [7:0] n10813_o;
  wire [7:0] n10814_o;
  wire [7:0] n10815_o;
  wire [7:0] n10816_o;
  wire [7:0] n10817_o;
  wire [7:0] n10818_o;
  wire [7:0] n10819_o;
  wire [7:0] n10820_o;
  wire [7:0] n10821_o;
  wire [7:0] n10822_o;
  wire [7:0] n10823_o;
  wire [7:0] n10824_o;
  wire [7:0] n10825_o;
  wire [7:0] n10826_o;
  wire [7:0] n10827_o;
  wire [7:0] n10828_o;
  wire [7:0] n10829_o;
  wire [7:0] n10830_o;
  wire [7:0] n10831_o;
  wire [7:0] n10832_o;
  wire [7:0] n10833_o;
  wire [7:0] n10834_o;
  wire [7:0] n10835_o;
  wire [7:0] n10836_o;
  wire [7:0] n10837_o;
  wire [7:0] n10838_o;
  wire [7:0] n10839_o;
  wire [7:0] n10840_o;
  wire [7:0] n10841_o;
  wire [7:0] n10842_o;
  wire [7:0] n10843_o;
  wire [7:0] n10844_o;
  wire [7:0] n10845_o;
  wire [7:0] n10846_o;
  wire [7:0] n10847_o;
  wire [7:0] n10848_o;
  wire [7:0] n10849_o;
  wire [7:0] n10850_o;
  wire [7:0] n10851_o;
  wire [7:0] n10852_o;
  wire [7:0] n10853_o;
  wire [7:0] n10854_o;
  wire [7:0] n10855_o;
  wire [7:0] n10856_o;
  wire [7:0] n10857_o;
  wire [7:0] n10858_o;
  wire [7:0] n10859_o;
  wire [7:0] n10860_o;
  wire [7:0] n10861_o;
  wire [7:0] n10862_o;
  wire [7:0] n10863_o;
  wire [7:0] n10864_o;
  wire [7:0] n10865_o;
  wire [7:0] n10866_o;
  wire [7:0] n10867_o;
  wire [7:0] n10868_o;
  wire [7:0] n10869_o;
  wire [7:0] n10870_o;
  wire [7:0] n10871_o;
  wire [7:0] n10872_o;
  wire [7:0] n10873_o;
  wire [7:0] n10874_o;
  wire [7:0] n10875_o;
  wire [7:0] n10876_o;
  wire [7:0] n10877_o;
  wire [7:0] n10878_o;
  wire [7:0] n10879_o;
  wire [7:0] n10880_o;
  wire [7:0] n10881_o;
  wire [7:0] n10882_o;
  wire [7:0] n10883_o;
  wire [7:0] n10884_o;
  wire [7:0] n10885_o;
  wire [7:0] n10886_o;
  wire [7:0] n10887_o;
  wire [7:0] n10888_o;
  wire [7:0] n10889_o;
  wire [7:0] n10890_o;
  wire [7:0] n10891_o;
  wire [7:0] n10892_o;
  wire [7:0] n10893_o;
  wire [7:0] n10894_o;
  wire [7:0] n10895_o;
  wire [7:0] n10896_o;
  wire [7:0] n10897_o;
  wire [7:0] n10898_o;
  wire [7:0] n10899_o;
  wire [7:0] n10900_o;
  wire [7:0] n10901_o;
  wire [7:0] n10902_o;
  wire [7:0] n10903_o;
  wire [7:0] n10904_o;
  wire [7:0] n10905_o;
  wire [7:0] n10906_o;
  wire [7:0] n10907_o;
  wire [7:0] n10908_o;
  wire [7:0] n10909_o;
  wire [7:0] n10910_o;
  wire [7:0] n10911_o;
  wire [7:0] n10912_o;
  wire [7:0] n10913_o;
  wire [7:0] n10914_o;
  wire [7:0] n10915_o;
  wire [7:0] n10916_o;
  wire [7:0] n10917_o;
  wire [7:0] n10918_o;
  wire [7:0] n10919_o;
  wire [7:0] n10920_o;
  wire [7:0] n10921_o;
  wire [7:0] n10922_o;
  wire [7:0] n10923_o;
  wire [7:0] n10924_o;
  wire [7:0] n10925_o;
  wire [7:0] n10926_o;
  wire [7:0] n10927_o;
  wire [7:0] n10928_o;
  wire [7:0] n10929_o;
  wire [7:0] n10930_o;
  wire [7:0] n10931_o;
  wire [7:0] n10932_o;
  wire [7:0] n10933_o;
  wire [7:0] n10934_o;
  wire [7:0] n10935_o;
  wire [7:0] n10936_o;
  wire [7:0] n10937_o;
  wire [7:0] n10938_o;
  wire [7:0] n10939_o;
  wire [7:0] n10940_o;
  wire [7:0] n10941_o;
  wire [7:0] n10942_o;
  wire [7:0] n10943_o;
  wire [7:0] n10944_o;
  wire [7:0] n10945_o;
  wire [7:0] n10946_o;
  wire [7:0] n10947_o;
  wire [7:0] n10948_o;
  wire [7:0] n10949_o;
  wire [7:0] n10950_o;
  wire [7:0] n10951_o;
  wire [7:0] n10952_o;
  wire [7:0] n10953_o;
  wire [7:0] n10954_o;
  wire [7:0] n10955_o;
  wire [7:0] n10956_o;
  wire [7:0] n10957_o;
  wire [7:0] n10958_o;
  wire [7:0] n10959_o;
  wire [7:0] n10960_o;
  wire [7:0] n10961_o;
  wire [7:0] n10962_o;
  wire [7:0] n10963_o;
  wire [7:0] n10964_o;
  wire [7:0] n10965_o;
  wire [7:0] n10966_o;
  wire [7:0] n10967_o;
  wire [7:0] n10968_o;
  wire [7:0] n10969_o;
  wire [7:0] n10970_o;
  wire [7:0] n10971_o;
  wire [7:0] n10972_o;
  wire [7:0] n10973_o;
  wire [7:0] n10974_o;
  wire [7:0] n10975_o;
  wire [7:0] n10976_o;
  wire [7:0] n10977_o;
  wire [7:0] n10978_o;
  wire [7:0] n10979_o;
  wire [7:0] n10980_o;
  wire [7:0] n10981_o;
  wire [7:0] n10982_o;
  wire [7:0] n10983_o;
  wire [7:0] n10984_o;
  wire [7:0] n10985_o;
  wire [7:0] n10986_o;
  wire [7:0] n10987_o;
  wire [7:0] n10988_o;
  wire [7:0] n10989_o;
  wire [7:0] n10990_o;
  wire [7:0] n10991_o;
  wire [7:0] n10992_o;
  wire [7:0] n10993_o;
  wire [7:0] n10994_o;
  wire [7:0] n10995_o;
  wire [7:0] n10996_o;
  wire [7:0] n10997_o;
  wire [7:0] n10998_o;
  wire [7:0] n10999_o;
  wire [7:0] n11000_o;
  wire [7:0] n11001_o;
  wire [7:0] n11002_o;
  wire [7:0] n11003_o;
  wire [7:0] n11004_o;
  wire [7:0] n11005_o;
  wire [7:0] n11006_o;
  wire [7:0] n11007_o;
  wire [7:0] n11008_o;
  wire [7:0] n11009_o;
  wire [7:0] n11010_o;
  wire [7:0] n11011_o;
  wire [7:0] n11012_o;
  wire [7:0] n11013_o;
  wire [7:0] n11014_o;
  wire [7:0] n11015_o;
  wire [7:0] n11016_o;
  wire [7:0] n11017_o;
  wire [7:0] n11018_o;
  wire [7:0] n11019_o;
  wire [7:0] n11020_o;
  wire [7:0] n11021_o;
  wire [7:0] n11022_o;
  wire [7:0] n11023_o;
  wire [7:0] n11024_o;
  wire [7:0] n11025_o;
  wire [7:0] n11026_o;
  wire [7:0] n11027_o;
  wire [7:0] n11028_o;
  wire [7:0] n11029_o;
  wire [7:0] n11030_o;
  wire [7:0] n11031_o;
  wire [7:0] n11032_o;
  wire [7:0] n11033_o;
  wire [7:0] n11034_o;
  wire [7:0] n11035_o;
  wire [7:0] n11036_o;
  wire [7:0] n11037_o;
  wire [7:0] n11038_o;
  wire [7:0] n11039_o;
  wire [7:0] n11040_o;
  wire [7:0] n11041_o;
  wire [7:0] n11042_o;
  wire [7:0] n11043_o;
  wire [7:0] n11044_o;
  wire [7:0] n11045_o;
  wire [7:0] n11046_o;
  wire [7:0] n11047_o;
  wire [7:0] n11048_o;
  wire [7:0] n11049_o;
  wire [7:0] n11050_o;
  wire [7:0] n11051_o;
  wire [7:0] n11052_o;
  wire [7:0] n11053_o;
  wire [7:0] n11054_o;
  wire [1:0] n11055_o;
  reg [7:0] n11056_o;
  wire [1:0] n11057_o;
  reg [7:0] n11058_o;
  wire [1:0] n11059_o;
  reg [7:0] n11060_o;
  wire [1:0] n11061_o;
  reg [7:0] n11062_o;
  wire [1:0] n11063_o;
  reg [7:0] n11064_o;
  wire [1:0] n11065_o;
  reg [7:0] n11066_o;
  wire [1:0] n11067_o;
  reg [7:0] n11068_o;
  wire [1:0] n11069_o;
  reg [7:0] n11070_o;
  wire [1:0] n11071_o;
  reg [7:0] n11072_o;
  wire [1:0] n11073_o;
  reg [7:0] n11074_o;
  wire [1:0] n11075_o;
  reg [7:0] n11076_o;
  wire [1:0] n11077_o;
  reg [7:0] n11078_o;
  wire [1:0] n11079_o;
  reg [7:0] n11080_o;
  wire [1:0] n11081_o;
  reg [7:0] n11082_o;
  wire [1:0] n11083_o;
  reg [7:0] n11084_o;
  wire [1:0] n11085_o;
  reg [7:0] n11086_o;
  wire [1:0] n11087_o;
  reg [7:0] n11088_o;
  wire [1:0] n11089_o;
  reg [7:0] n11090_o;
  wire [1:0] n11091_o;
  reg [7:0] n11092_o;
  wire [1:0] n11093_o;
  reg [7:0] n11094_o;
  wire [1:0] n11095_o;
  reg [7:0] n11096_o;
  wire [1:0] n11097_o;
  reg [7:0] n11098_o;
  wire [1:0] n11099_o;
  reg [7:0] n11100_o;
  wire [1:0] n11101_o;
  reg [7:0] n11102_o;
  wire [1:0] n11103_o;
  reg [7:0] n11104_o;
  wire [1:0] n11105_o;
  reg [7:0] n11106_o;
  wire [1:0] n11107_o;
  reg [7:0] n11108_o;
  wire [1:0] n11109_o;
  reg [7:0] n11110_o;
  wire [1:0] n11111_o;
  reg [7:0] n11112_o;
  wire [1:0] n11113_o;
  reg [7:0] n11114_o;
  wire [1:0] n11115_o;
  reg [7:0] n11116_o;
  wire [1:0] n11117_o;
  reg [7:0] n11118_o;
  wire [1:0] n11119_o;
  reg [7:0] n11120_o;
  wire [1:0] n11121_o;
  reg [7:0] n11122_o;
  wire [1:0] n11123_o;
  reg [7:0] n11124_o;
  wire [1:0] n11125_o;
  reg [7:0] n11126_o;
  wire [1:0] n11127_o;
  reg [7:0] n11128_o;
  wire [1:0] n11129_o;
  reg [7:0] n11130_o;
  wire [1:0] n11131_o;
  reg [7:0] n11132_o;
  wire [1:0] n11133_o;
  reg [7:0] n11134_o;
  wire [1:0] n11135_o;
  reg [7:0] n11136_o;
  wire [1:0] n11137_o;
  reg [7:0] n11138_o;
  wire [1:0] n11139_o;
  reg [7:0] n11140_o;
  wire [1:0] n11141_o;
  reg [7:0] n11142_o;
  wire [1:0] n11143_o;
  reg [7:0] n11144_o;
  wire [1:0] n11145_o;
  reg [7:0] n11146_o;
  wire [1:0] n11147_o;
  reg [7:0] n11148_o;
  wire [1:0] n11149_o;
  reg [7:0] n11150_o;
  wire [1:0] n11151_o;
  reg [7:0] n11152_o;
  wire [1:0] n11153_o;
  reg [7:0] n11154_o;
  wire [1:0] n11155_o;
  reg [7:0] n11156_o;
  wire [1:0] n11157_o;
  reg [7:0] n11158_o;
  wire [1:0] n11159_o;
  reg [7:0] n11160_o;
  wire [1:0] n11161_o;
  reg [7:0] n11162_o;
  wire [1:0] n11163_o;
  reg [7:0] n11164_o;
  wire [1:0] n11165_o;
  reg [7:0] n11166_o;
  wire [1:0] n11167_o;
  reg [7:0] n11168_o;
  wire [1:0] n11169_o;
  reg [7:0] n11170_o;
  wire [1:0] n11171_o;
  reg [7:0] n11172_o;
  wire [1:0] n11173_o;
  reg [7:0] n11174_o;
  wire [1:0] n11175_o;
  reg [7:0] n11176_o;
  wire [1:0] n11177_o;
  reg [7:0] n11178_o;
  wire [1:0] n11179_o;
  reg [7:0] n11180_o;
  wire [1:0] n11181_o;
  reg [7:0] n11182_o;
  wire [1:0] n11183_o;
  reg [7:0] n11184_o;
  wire [1:0] n11185_o;
  reg [7:0] n11186_o;
  wire [1:0] n11187_o;
  reg [7:0] n11188_o;
  wire [1:0] n11189_o;
  reg [7:0] n11190_o;
  wire [1:0] n11191_o;
  reg [7:0] n11192_o;
  wire [1:0] n11193_o;
  reg [7:0] n11194_o;
  wire [1:0] n11195_o;
  reg [7:0] n11196_o;
  wire [1:0] n11197_o;
  reg [7:0] n11198_o;
  wire [1:0] n11199_o;
  reg [7:0] n11200_o;
  wire [1:0] n11201_o;
  reg [7:0] n11202_o;
  wire [1:0] n11203_o;
  reg [7:0] n11204_o;
  wire [1:0] n11205_o;
  reg [7:0] n11206_o;
  wire [1:0] n11207_o;
  reg [7:0] n11208_o;
  wire [1:0] n11209_o;
  reg [7:0] n11210_o;
  wire [1:0] n11211_o;
  reg [7:0] n11212_o;
  wire [1:0] n11213_o;
  reg [7:0] n11214_o;
  wire [1:0] n11215_o;
  reg [7:0] n11216_o;
  wire [1:0] n11217_o;
  reg [7:0] n11218_o;
  wire [1:0] n11219_o;
  reg [7:0] n11220_o;
  wire [1:0] n11221_o;
  reg [7:0] n11222_o;
  wire [1:0] n11223_o;
  reg [7:0] n11224_o;
  assign half_o = n9758_q;
  assign free_o = n9759_q;
  assign rdata_o = n9760_q;
  assign avail_o = n9761_q;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:84:10  */
  assign fifo = n9757_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:87:10  */
  assign level_diff = n9703_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:99:19  */
  assign n9645_o = 1'b0 ? re_i : n9647_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:99:64  */
  assign n9646_o = fifo[2081];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:99:55  */
  assign n9647_o = re_i & n9646_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:100:19  */
  assign n9649_o = 1'b0 ? we_i : n9651_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:100:64  */
  assign n9650_o = fifo[2080];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:100:55  */
  assign n9651_o = we_i & n9650_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:107:16  */
  assign n9653_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:114:19  */
  assign n9658_o = fifo[0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:115:55  */
  assign n9659_o = fifo[10:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:115:62  */
  assign n9661_o = n9659_o + 9'b000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:519:52  */
  assign n9662_o = fifo[10:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:114:7  */
  assign n9663_o = n9658_o ? n9661_o : n9662_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:112:7  */
  assign n9664_o = clear_i ? 9'b000000000 : n9663_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:120:19  */
  assign n9666_o = fifo[1];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:121:55  */
  assign n9667_o = fifo[19:11];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:121:62  */
  assign n9669_o = n9667_o + 9'b000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:266:16  */
  assign n9670_o = fifo[19:11];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:120:7  */
  assign n9671_o = n9666_o ? n9669_o : n9670_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:118:7  */
  assign n9672_o = clear_i ? 9'b000000000 : n9671_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:177:7  */
  assign n9673_o = {n9672_o, n9664_o};
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:186:27  */
  assign n9676_o = {9'b000000000, 9'b000000000};
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:131:39  */
  assign n9680_o = fifo[18:11];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:131:80  */
  assign n9681_o = fifo[9:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:131:68  */
  assign n9682_o = n9680_o == n9681_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:131:23  */
  assign n9683_o = n9682_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:132:39  */
  assign n9686_o = fifo[19];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:132:70  */
  assign n9687_o = fifo[10];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:132:57  */
  assign n9688_o = n9686_o != n9687_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:132:99  */
  assign n9689_o = fifo[2076];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:132:89  */
  assign n9690_o = n9688_o & n9689_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:132:23  */
  assign n9691_o = n9690_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:133:39  */
  assign n9694_o = fifo[19];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:133:70  */
  assign n9695_o = fifo[10];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:133:58  */
  assign n9696_o = n9694_o == n9695_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:133:99  */
  assign n9697_o = fifo[2076];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:133:89  */
  assign n9698_o = n9696_o & n9697_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:133:23  */
  assign n9699_o = n9698_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:134:51  */
  assign n9701_o = fifo[10:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:134:74  */
  assign n9702_o = fifo[19:11];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:134:58  */
  assign n9703_o = n9701_o - n9702_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:135:29  */
  assign n9704_o = level_diff[7];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:135:57  */
  assign n9705_o = fifo[2078];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:135:49  */
  assign n9706_o = n9704_o | n9705_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:146:26  */
  assign n9707_o = fifo[2078];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:146:17  */
  assign n9708_o = ~n9707_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:147:26  */
  assign n9709_o = fifo[2077];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:147:17  */
  assign n9710_o = ~n9709_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:163:18  */
  assign n9712_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:168:25  */
  assign n9714_o = fifo[2080];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:169:25  */
  assign n9715_o = fifo[2081];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:170:25  */
  assign n9716_o = fifo[2079];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:183:18  */
  assign n9729_o = fifo[0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:51  */
  assign n9730_o = fifo[9:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:21  */
  assign n9733_o = 8'b11111111 - n9730_o;
  assign n9735_o = fifo[2067:20];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:62  */
  assign n9745_o = fifo[18:11];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:32  */
  assign n9748_o = 8'b11111111 - n9745_o;
  assign n9753_o = fifo[2067:20];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:182:7  */
  assign n9754_o = n9729_o ? n10798_o : n9753_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:182:7  */
  always @(posedge clk_i)
    n9755_q <= n9754_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:110:5  */
  always @(posedge clk_i or posedge n9653_o)
    if (n9653_o)
      n9756_q <= n9676_o;
    else
      n9756_q <= n9673_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:107:5  */
  assign n9757_o = {n9710_o, n9708_o, n9706_o, n9691_o, n9699_o, n9683_o, 8'b00000000, n9755_q, n9756_q, n9645_o, n9649_o};
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:167:7  */
  always @(posedge clk_i or posedge n9712_o)
    if (n9712_o)
      n9758_q <= 1'b0;
    else
      n9758_q <= n9716_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:167:7  */
  always @(posedge clk_i or posedge n9712_o)
    if (n9712_o)
      n9759_q <= 1'b0;
    else
      n9759_q <= n9714_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:223:7  */
  always @(posedge clk_i)
    n9760_q <= n11224_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:167:7  */
  always @(posedge clk_i or posedge n9712_o)
    if (n9712_o)
      n9761_q <= 1'b0;
    else
      n9761_q <= n9715_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9762_o = n9733_o[7];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9763_o = ~n9762_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9764_o = n9733_o[6];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9765_o = ~n9764_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9766_o = n9763_o & n9765_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9767_o = n9763_o & n9764_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9768_o = n9762_o & n9765_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9769_o = n9762_o & n9764_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9770_o = n9733_o[5];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9771_o = ~n9770_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9772_o = n9766_o & n9771_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9773_o = n9766_o & n9770_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9774_o = n9767_o & n9771_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9775_o = n9767_o & n9770_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9776_o = n9768_o & n9771_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9777_o = n9768_o & n9770_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9778_o = n9769_o & n9771_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9779_o = n9769_o & n9770_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9780_o = n9733_o[4];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9781_o = ~n9780_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9782_o = n9772_o & n9781_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9783_o = n9772_o & n9780_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9784_o = n9773_o & n9781_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9785_o = n9773_o & n9780_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9786_o = n9774_o & n9781_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9787_o = n9774_o & n9780_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9788_o = n9775_o & n9781_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9789_o = n9775_o & n9780_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9790_o = n9776_o & n9781_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9791_o = n9776_o & n9780_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9792_o = n9777_o & n9781_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9793_o = n9777_o & n9780_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9794_o = n9778_o & n9781_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9795_o = n9778_o & n9780_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9796_o = n9779_o & n9781_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9797_o = n9779_o & n9780_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9798_o = n9733_o[3];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9799_o = ~n9798_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9800_o = n9782_o & n9799_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9801_o = n9782_o & n9798_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9802_o = n9783_o & n9799_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9803_o = n9783_o & n9798_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9804_o = n9784_o & n9799_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9805_o = n9784_o & n9798_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9806_o = n9785_o & n9799_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9807_o = n9785_o & n9798_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9808_o = n9786_o & n9799_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9809_o = n9786_o & n9798_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9810_o = n9787_o & n9799_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9811_o = n9787_o & n9798_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9812_o = n9788_o & n9799_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9813_o = n9788_o & n9798_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9814_o = n9789_o & n9799_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9815_o = n9789_o & n9798_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9816_o = n9790_o & n9799_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9817_o = n9790_o & n9798_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9818_o = n9791_o & n9799_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9819_o = n9791_o & n9798_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9820_o = n9792_o & n9799_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9821_o = n9792_o & n9798_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9822_o = n9793_o & n9799_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9823_o = n9793_o & n9798_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9824_o = n9794_o & n9799_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9825_o = n9794_o & n9798_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9826_o = n9795_o & n9799_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9827_o = n9795_o & n9798_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9828_o = n9796_o & n9799_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9829_o = n9796_o & n9798_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9830_o = n9797_o & n9799_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9831_o = n9797_o & n9798_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9832_o = n9733_o[2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9833_o = ~n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9834_o = n9800_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9835_o = n9800_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9836_o = n9801_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9837_o = n9801_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9838_o = n9802_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9839_o = n9802_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9840_o = n9803_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9841_o = n9803_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9842_o = n9804_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9843_o = n9804_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9844_o = n9805_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9845_o = n9805_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9846_o = n9806_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9847_o = n9806_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9848_o = n9807_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9849_o = n9807_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9850_o = n9808_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9851_o = n9808_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9852_o = n9809_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9853_o = n9809_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9854_o = n9810_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9855_o = n9810_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9856_o = n9811_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9857_o = n9811_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9858_o = n9812_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9859_o = n9812_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9860_o = n9813_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9861_o = n9813_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9862_o = n9814_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9863_o = n9814_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9864_o = n9815_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9865_o = n9815_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9866_o = n9816_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9867_o = n9816_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9868_o = n9817_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9869_o = n9817_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9870_o = n9818_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9871_o = n9818_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9872_o = n9819_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9873_o = n9819_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9874_o = n9820_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9875_o = n9820_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9876_o = n9821_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9877_o = n9821_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9878_o = n9822_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9879_o = n9822_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9880_o = n9823_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9881_o = n9823_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9882_o = n9824_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9883_o = n9824_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9884_o = n9825_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9885_o = n9825_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9886_o = n9826_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9887_o = n9826_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9888_o = n9827_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9889_o = n9827_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9890_o = n9828_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9891_o = n9828_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9892_o = n9829_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9893_o = n9829_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9894_o = n9830_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9895_o = n9830_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9896_o = n9831_o & n9833_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9897_o = n9831_o & n9832_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9898_o = n9733_o[1];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9899_o = ~n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9900_o = n9834_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9901_o = n9834_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9902_o = n9835_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9903_o = n9835_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9904_o = n9836_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9905_o = n9836_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9906_o = n9837_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9907_o = n9837_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9908_o = n9838_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9909_o = n9838_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9910_o = n9839_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9911_o = n9839_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9912_o = n9840_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9913_o = n9840_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9914_o = n9841_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9915_o = n9841_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9916_o = n9842_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9917_o = n9842_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9918_o = n9843_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9919_o = n9843_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9920_o = n9844_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9921_o = n9844_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9922_o = n9845_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9923_o = n9845_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9924_o = n9846_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9925_o = n9846_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9926_o = n9847_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9927_o = n9847_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9928_o = n9848_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9929_o = n9848_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9930_o = n9849_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9931_o = n9849_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9932_o = n9850_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9933_o = n9850_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9934_o = n9851_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9935_o = n9851_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9936_o = n9852_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9937_o = n9852_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9938_o = n9853_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9939_o = n9853_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9940_o = n9854_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9941_o = n9854_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9942_o = n9855_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9943_o = n9855_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9944_o = n9856_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9945_o = n9856_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9946_o = n9857_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9947_o = n9857_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9948_o = n9858_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9949_o = n9858_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9950_o = n9859_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9951_o = n9859_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9952_o = n9860_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9953_o = n9860_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9954_o = n9861_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9955_o = n9861_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9956_o = n9862_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9957_o = n9862_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9958_o = n9863_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9959_o = n9863_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9960_o = n9864_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9961_o = n9864_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9962_o = n9865_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9963_o = n9865_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9964_o = n9866_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9965_o = n9866_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9966_o = n9867_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9967_o = n9867_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9968_o = n9868_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9969_o = n9868_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9970_o = n9869_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9971_o = n9869_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9972_o = n9870_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9973_o = n9870_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9974_o = n9871_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9975_o = n9871_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9976_o = n9872_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9977_o = n9872_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9978_o = n9873_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9979_o = n9873_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9980_o = n9874_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9981_o = n9874_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9982_o = n9875_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9983_o = n9875_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9984_o = n9876_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9985_o = n9876_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9986_o = n9877_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9987_o = n9877_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9988_o = n9878_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9989_o = n9878_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9990_o = n9879_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9991_o = n9879_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9992_o = n9880_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9993_o = n9880_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9994_o = n9881_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9995_o = n9881_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9996_o = n9882_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9997_o = n9882_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9998_o = n9883_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n9999_o = n9883_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10000_o = n9884_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10001_o = n9884_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10002_o = n9885_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10003_o = n9885_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10004_o = n9886_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10005_o = n9886_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10006_o = n9887_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10007_o = n9887_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10008_o = n9888_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10009_o = n9888_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10010_o = n9889_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10011_o = n9889_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10012_o = n9890_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10013_o = n9890_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10014_o = n9891_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10015_o = n9891_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10016_o = n9892_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10017_o = n9892_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10018_o = n9893_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10019_o = n9893_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10020_o = n9894_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10021_o = n9894_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10022_o = n9895_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10023_o = n9895_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10024_o = n9896_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10025_o = n9896_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10026_o = n9897_o & n9899_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10027_o = n9897_o & n9898_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10028_o = n9733_o[0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10029_o = ~n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10030_o = n9900_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10031_o = n9900_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10032_o = n9901_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10033_o = n9901_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10034_o = n9902_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10035_o = n9902_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10036_o = n9903_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10037_o = n9903_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10038_o = n9904_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10039_o = n9904_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10040_o = n9905_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10041_o = n9905_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10042_o = n9906_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10043_o = n9906_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10044_o = n9907_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10045_o = n9907_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10046_o = n9908_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10047_o = n9908_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10048_o = n9909_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10049_o = n9909_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10050_o = n9910_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10051_o = n9910_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10052_o = n9911_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10053_o = n9911_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10054_o = n9912_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10055_o = n9912_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10056_o = n9913_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10057_o = n9913_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10058_o = n9914_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10059_o = n9914_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10060_o = n9915_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10061_o = n9915_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10062_o = n9916_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10063_o = n9916_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10064_o = n9917_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10065_o = n9917_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10066_o = n9918_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10067_o = n9918_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10068_o = n9919_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10069_o = n9919_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10070_o = n9920_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10071_o = n9920_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10072_o = n9921_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10073_o = n9921_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10074_o = n9922_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10075_o = n9922_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10076_o = n9923_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10077_o = n9923_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10078_o = n9924_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10079_o = n9924_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10080_o = n9925_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10081_o = n9925_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10082_o = n9926_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10083_o = n9926_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10084_o = n9927_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10085_o = n9927_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10086_o = n9928_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10087_o = n9928_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10088_o = n9929_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10089_o = n9929_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10090_o = n9930_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10091_o = n9930_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10092_o = n9931_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10093_o = n9931_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10094_o = n9932_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10095_o = n9932_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10096_o = n9933_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10097_o = n9933_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10098_o = n9934_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10099_o = n9934_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10100_o = n9935_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10101_o = n9935_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10102_o = n9936_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10103_o = n9936_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10104_o = n9937_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10105_o = n9937_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10106_o = n9938_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10107_o = n9938_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10108_o = n9939_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10109_o = n9939_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10110_o = n9940_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10111_o = n9940_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10112_o = n9941_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10113_o = n9941_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10114_o = n9942_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10115_o = n9942_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10116_o = n9943_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10117_o = n9943_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10118_o = n9944_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10119_o = n9944_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10120_o = n9945_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10121_o = n9945_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10122_o = n9946_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10123_o = n9946_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10124_o = n9947_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10125_o = n9947_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10126_o = n9948_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10127_o = n9948_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10128_o = n9949_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10129_o = n9949_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10130_o = n9950_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10131_o = n9950_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10132_o = n9951_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10133_o = n9951_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10134_o = n9952_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10135_o = n9952_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10136_o = n9953_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10137_o = n9953_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10138_o = n9954_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10139_o = n9954_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10140_o = n9955_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10141_o = n9955_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10142_o = n9956_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10143_o = n9956_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10144_o = n9957_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10145_o = n9957_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10146_o = n9958_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10147_o = n9958_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10148_o = n9959_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10149_o = n9959_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10150_o = n9960_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10151_o = n9960_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10152_o = n9961_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10153_o = n9961_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10154_o = n9962_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10155_o = n9962_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10156_o = n9963_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10157_o = n9963_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10158_o = n9964_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10159_o = n9964_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10160_o = n9965_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10161_o = n9965_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10162_o = n9966_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10163_o = n9966_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10164_o = n9967_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10165_o = n9967_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10166_o = n9968_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10167_o = n9968_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10168_o = n9969_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10169_o = n9969_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10170_o = n9970_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10171_o = n9970_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10172_o = n9971_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10173_o = n9971_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10174_o = n9972_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10175_o = n9972_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10176_o = n9973_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10177_o = n9973_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10178_o = n9974_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10179_o = n9974_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10180_o = n9975_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10181_o = n9975_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10182_o = n9976_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10183_o = n9976_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10184_o = n9977_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10185_o = n9977_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10186_o = n9978_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10187_o = n9978_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10188_o = n9979_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10189_o = n9979_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10190_o = n9980_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10191_o = n9980_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10192_o = n9981_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10193_o = n9981_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10194_o = n9982_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10195_o = n9982_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10196_o = n9983_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10197_o = n9983_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10198_o = n9984_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10199_o = n9984_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10200_o = n9985_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10201_o = n9985_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10202_o = n9986_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10203_o = n9986_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10204_o = n9987_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10205_o = n9987_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10206_o = n9988_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10207_o = n9988_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10208_o = n9989_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10209_o = n9989_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10210_o = n9990_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10211_o = n9990_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10212_o = n9991_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10213_o = n9991_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10214_o = n9992_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10215_o = n9992_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10216_o = n9993_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10217_o = n9993_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10218_o = n9994_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10219_o = n9994_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10220_o = n9995_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10221_o = n9995_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10222_o = n9996_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10223_o = n9996_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10224_o = n9997_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10225_o = n9997_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10226_o = n9998_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10227_o = n9998_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10228_o = n9999_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10229_o = n9999_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10230_o = n10000_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10231_o = n10000_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10232_o = n10001_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10233_o = n10001_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10234_o = n10002_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10235_o = n10002_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10236_o = n10003_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10237_o = n10003_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10238_o = n10004_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10239_o = n10004_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10240_o = n10005_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10241_o = n10005_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10242_o = n10006_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10243_o = n10006_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10244_o = n10007_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10245_o = n10007_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10246_o = n10008_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10247_o = n10008_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10248_o = n10009_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10249_o = n10009_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10250_o = n10010_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10251_o = n10010_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10252_o = n10011_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10253_o = n10011_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10254_o = n10012_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10255_o = n10012_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10256_o = n10013_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10257_o = n10013_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10258_o = n10014_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10259_o = n10014_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10260_o = n10015_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10261_o = n10015_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10262_o = n10016_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10263_o = n10016_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10264_o = n10017_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10265_o = n10017_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10266_o = n10018_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10267_o = n10018_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10268_o = n10019_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10269_o = n10019_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10270_o = n10020_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10271_o = n10020_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10272_o = n10021_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10273_o = n10021_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10274_o = n10022_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10275_o = n10022_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10276_o = n10023_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10277_o = n10023_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10278_o = n10024_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10279_o = n10024_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10280_o = n10025_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10281_o = n10025_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10282_o = n10026_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10283_o = n10026_o & n10028_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10284_o = n10027_o & n10029_o;
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10285_o = n10027_o & n10028_o;
  assign n10286_o = n9735_o[7:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10287_o = n10030_o ? wdata_i : n10286_o;
  assign n10288_o = n9735_o[15:8];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10289_o = n10031_o ? wdata_i : n10288_o;
  assign n10290_o = n9735_o[23:16];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10291_o = n10032_o ? wdata_i : n10290_o;
  assign n10292_o = n9735_o[31:24];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10293_o = n10033_o ? wdata_i : n10292_o;
  assign n10294_o = n9735_o[39:32];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10295_o = n10034_o ? wdata_i : n10294_o;
  assign n10296_o = n9735_o[47:40];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10297_o = n10035_o ? wdata_i : n10296_o;
  assign n10298_o = n9735_o[55:48];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10299_o = n10036_o ? wdata_i : n10298_o;
  assign n10300_o = n9735_o[63:56];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10301_o = n10037_o ? wdata_i : n10300_o;
  assign n10302_o = n9735_o[71:64];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10303_o = n10038_o ? wdata_i : n10302_o;
  assign n10304_o = n9735_o[79:72];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10305_o = n10039_o ? wdata_i : n10304_o;
  assign n10306_o = n9735_o[87:80];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10307_o = n10040_o ? wdata_i : n10306_o;
  assign n10308_o = n9735_o[95:88];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10309_o = n10041_o ? wdata_i : n10308_o;
  assign n10310_o = n9735_o[103:96];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10311_o = n10042_o ? wdata_i : n10310_o;
  assign n10312_o = n9735_o[111:104];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10313_o = n10043_o ? wdata_i : n10312_o;
  assign n10314_o = n9735_o[119:112];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10315_o = n10044_o ? wdata_i : n10314_o;
  assign n10316_o = n9735_o[127:120];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10317_o = n10045_o ? wdata_i : n10316_o;
  assign n10318_o = n9735_o[135:128];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10319_o = n10046_o ? wdata_i : n10318_o;
  assign n10320_o = n9735_o[143:136];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10321_o = n10047_o ? wdata_i : n10320_o;
  assign n10322_o = n9735_o[151:144];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10323_o = n10048_o ? wdata_i : n10322_o;
  assign n10324_o = n9735_o[159:152];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10325_o = n10049_o ? wdata_i : n10324_o;
  assign n10326_o = n9735_o[167:160];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10327_o = n10050_o ? wdata_i : n10326_o;
  assign n10328_o = n9735_o[175:168];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10329_o = n10051_o ? wdata_i : n10328_o;
  assign n10330_o = n9735_o[183:176];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10331_o = n10052_o ? wdata_i : n10330_o;
  assign n10332_o = n9735_o[191:184];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10333_o = n10053_o ? wdata_i : n10332_o;
  assign n10334_o = n9735_o[199:192];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10335_o = n10054_o ? wdata_i : n10334_o;
  assign n10336_o = n9735_o[207:200];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10337_o = n10055_o ? wdata_i : n10336_o;
  assign n10338_o = n9735_o[215:208];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10339_o = n10056_o ? wdata_i : n10338_o;
  assign n10340_o = n9735_o[223:216];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10341_o = n10057_o ? wdata_i : n10340_o;
  assign n10342_o = n9735_o[231:224];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10343_o = n10058_o ? wdata_i : n10342_o;
  assign n10344_o = n9735_o[239:232];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10345_o = n10059_o ? wdata_i : n10344_o;
  assign n10346_o = n9735_o[247:240];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10347_o = n10060_o ? wdata_i : n10346_o;
  assign n10348_o = n9735_o[255:248];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10349_o = n10061_o ? wdata_i : n10348_o;
  assign n10350_o = n9735_o[263:256];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10351_o = n10062_o ? wdata_i : n10350_o;
  assign n10352_o = n9735_o[271:264];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10353_o = n10063_o ? wdata_i : n10352_o;
  assign n10354_o = n9735_o[279:272];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10355_o = n10064_o ? wdata_i : n10354_o;
  assign n10356_o = n9735_o[287:280];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10357_o = n10065_o ? wdata_i : n10356_o;
  assign n10358_o = n9735_o[295:288];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10359_o = n10066_o ? wdata_i : n10358_o;
  assign n10360_o = n9735_o[303:296];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10361_o = n10067_o ? wdata_i : n10360_o;
  assign n10362_o = n9735_o[311:304];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10363_o = n10068_o ? wdata_i : n10362_o;
  assign n10364_o = n9735_o[319:312];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10365_o = n10069_o ? wdata_i : n10364_o;
  assign n10366_o = n9735_o[327:320];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10367_o = n10070_o ? wdata_i : n10366_o;
  assign n10368_o = n9735_o[335:328];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10369_o = n10071_o ? wdata_i : n10368_o;
  assign n10370_o = n9735_o[343:336];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10371_o = n10072_o ? wdata_i : n10370_o;
  assign n10372_o = n9735_o[351:344];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10373_o = n10073_o ? wdata_i : n10372_o;
  assign n10374_o = n9735_o[359:352];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10375_o = n10074_o ? wdata_i : n10374_o;
  assign n10376_o = n9735_o[367:360];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10377_o = n10075_o ? wdata_i : n10376_o;
  assign n10378_o = n9735_o[375:368];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10379_o = n10076_o ? wdata_i : n10378_o;
  assign n10380_o = n9735_o[383:376];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10381_o = n10077_o ? wdata_i : n10380_o;
  assign n10382_o = n9735_o[391:384];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10383_o = n10078_o ? wdata_i : n10382_o;
  assign n10384_o = n9735_o[399:392];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10385_o = n10079_o ? wdata_i : n10384_o;
  assign n10386_o = n9735_o[407:400];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10387_o = n10080_o ? wdata_i : n10386_o;
  assign n10388_o = n9735_o[415:408];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10389_o = n10081_o ? wdata_i : n10388_o;
  assign n10390_o = n9735_o[423:416];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10391_o = n10082_o ? wdata_i : n10390_o;
  assign n10392_o = n9735_o[431:424];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10393_o = n10083_o ? wdata_i : n10392_o;
  assign n10394_o = n9735_o[439:432];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10395_o = n10084_o ? wdata_i : n10394_o;
  assign n10396_o = n9735_o[447:440];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10397_o = n10085_o ? wdata_i : n10396_o;
  assign n10398_o = n9735_o[455:448];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10399_o = n10086_o ? wdata_i : n10398_o;
  assign n10400_o = n9735_o[463:456];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10401_o = n10087_o ? wdata_i : n10400_o;
  assign n10402_o = n9735_o[471:464];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10403_o = n10088_o ? wdata_i : n10402_o;
  assign n10404_o = n9735_o[479:472];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10405_o = n10089_o ? wdata_i : n10404_o;
  assign n10406_o = n9735_o[487:480];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10407_o = n10090_o ? wdata_i : n10406_o;
  assign n10408_o = n9735_o[495:488];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10409_o = n10091_o ? wdata_i : n10408_o;
  assign n10410_o = n9735_o[503:496];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10411_o = n10092_o ? wdata_i : n10410_o;
  assign n10412_o = n9735_o[511:504];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10413_o = n10093_o ? wdata_i : n10412_o;
  assign n10414_o = n9735_o[519:512];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10415_o = n10094_o ? wdata_i : n10414_o;
  assign n10416_o = n9735_o[527:520];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10417_o = n10095_o ? wdata_i : n10416_o;
  assign n10418_o = n9735_o[535:528];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10419_o = n10096_o ? wdata_i : n10418_o;
  assign n10420_o = n9735_o[543:536];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10421_o = n10097_o ? wdata_i : n10420_o;
  assign n10422_o = n9735_o[551:544];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10423_o = n10098_o ? wdata_i : n10422_o;
  assign n10424_o = n9735_o[559:552];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10425_o = n10099_o ? wdata_i : n10424_o;
  assign n10426_o = n9735_o[567:560];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10427_o = n10100_o ? wdata_i : n10426_o;
  assign n10428_o = n9735_o[575:568];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10429_o = n10101_o ? wdata_i : n10428_o;
  assign n10430_o = n9735_o[583:576];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10431_o = n10102_o ? wdata_i : n10430_o;
  assign n10432_o = n9735_o[591:584];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10433_o = n10103_o ? wdata_i : n10432_o;
  assign n10434_o = n9735_o[599:592];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10435_o = n10104_o ? wdata_i : n10434_o;
  assign n10436_o = n9735_o[607:600];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10437_o = n10105_o ? wdata_i : n10436_o;
  assign n10438_o = n9735_o[615:608];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10439_o = n10106_o ? wdata_i : n10438_o;
  assign n10440_o = n9735_o[623:616];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10441_o = n10107_o ? wdata_i : n10440_o;
  assign n10442_o = n9735_o[631:624];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10443_o = n10108_o ? wdata_i : n10442_o;
  assign n10444_o = n9735_o[639:632];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10445_o = n10109_o ? wdata_i : n10444_o;
  assign n10446_o = n9735_o[647:640];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10447_o = n10110_o ? wdata_i : n10446_o;
  assign n10448_o = n9735_o[655:648];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10449_o = n10111_o ? wdata_i : n10448_o;
  assign n10450_o = n9735_o[663:656];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10451_o = n10112_o ? wdata_i : n10450_o;
  assign n10452_o = n9735_o[671:664];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10453_o = n10113_o ? wdata_i : n10452_o;
  assign n10454_o = n9735_o[679:672];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10455_o = n10114_o ? wdata_i : n10454_o;
  assign n10456_o = n9735_o[687:680];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10457_o = n10115_o ? wdata_i : n10456_o;
  assign n10458_o = n9735_o[695:688];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10459_o = n10116_o ? wdata_i : n10458_o;
  assign n10460_o = n9735_o[703:696];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10461_o = n10117_o ? wdata_i : n10460_o;
  assign n10462_o = n9735_o[711:704];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10463_o = n10118_o ? wdata_i : n10462_o;
  assign n10464_o = n9735_o[719:712];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10465_o = n10119_o ? wdata_i : n10464_o;
  assign n10466_o = n9735_o[727:720];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10467_o = n10120_o ? wdata_i : n10466_o;
  assign n10468_o = n9735_o[735:728];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10469_o = n10121_o ? wdata_i : n10468_o;
  assign n10470_o = n9735_o[743:736];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10471_o = n10122_o ? wdata_i : n10470_o;
  assign n10472_o = n9735_o[751:744];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10473_o = n10123_o ? wdata_i : n10472_o;
  assign n10474_o = n9735_o[759:752];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10475_o = n10124_o ? wdata_i : n10474_o;
  assign n10476_o = n9735_o[767:760];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10477_o = n10125_o ? wdata_i : n10476_o;
  assign n10478_o = n9735_o[775:768];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10479_o = n10126_o ? wdata_i : n10478_o;
  assign n10480_o = n9735_o[783:776];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10481_o = n10127_o ? wdata_i : n10480_o;
  assign n10482_o = n9735_o[791:784];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10483_o = n10128_o ? wdata_i : n10482_o;
  assign n10484_o = n9735_o[799:792];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10485_o = n10129_o ? wdata_i : n10484_o;
  assign n10486_o = n9735_o[807:800];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10487_o = n10130_o ? wdata_i : n10486_o;
  assign n10488_o = n9735_o[815:808];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10489_o = n10131_o ? wdata_i : n10488_o;
  assign n10490_o = n9735_o[823:816];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10491_o = n10132_o ? wdata_i : n10490_o;
  assign n10492_o = n9735_o[831:824];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10493_o = n10133_o ? wdata_i : n10492_o;
  assign n10494_o = n9735_o[839:832];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10495_o = n10134_o ? wdata_i : n10494_o;
  assign n10496_o = n9735_o[847:840];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10497_o = n10135_o ? wdata_i : n10496_o;
  assign n10498_o = n9735_o[855:848];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10499_o = n10136_o ? wdata_i : n10498_o;
  assign n10500_o = n9735_o[863:856];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10501_o = n10137_o ? wdata_i : n10500_o;
  assign n10502_o = n9735_o[871:864];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10503_o = n10138_o ? wdata_i : n10502_o;
  assign n10504_o = n9735_o[879:872];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10505_o = n10139_o ? wdata_i : n10504_o;
  assign n10506_o = n9735_o[887:880];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10507_o = n10140_o ? wdata_i : n10506_o;
  assign n10508_o = n9735_o[895:888];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10509_o = n10141_o ? wdata_i : n10508_o;
  assign n10510_o = n9735_o[903:896];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10511_o = n10142_o ? wdata_i : n10510_o;
  assign n10512_o = n9735_o[911:904];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10513_o = n10143_o ? wdata_i : n10512_o;
  assign n10514_o = n9735_o[919:912];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10515_o = n10144_o ? wdata_i : n10514_o;
  assign n10516_o = n9735_o[927:920];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10517_o = n10145_o ? wdata_i : n10516_o;
  assign n10518_o = n9735_o[935:928];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10519_o = n10146_o ? wdata_i : n10518_o;
  assign n10520_o = n9735_o[943:936];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10521_o = n10147_o ? wdata_i : n10520_o;
  assign n10522_o = n9735_o[951:944];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10523_o = n10148_o ? wdata_i : n10522_o;
  assign n10524_o = n9735_o[959:952];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10525_o = n10149_o ? wdata_i : n10524_o;
  assign n10526_o = n9735_o[967:960];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10527_o = n10150_o ? wdata_i : n10526_o;
  assign n10528_o = n9735_o[975:968];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10529_o = n10151_o ? wdata_i : n10528_o;
  assign n10530_o = n9735_o[983:976];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10531_o = n10152_o ? wdata_i : n10530_o;
  assign n10532_o = n9735_o[991:984];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10533_o = n10153_o ? wdata_i : n10532_o;
  assign n10534_o = n9735_o[999:992];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10535_o = n10154_o ? wdata_i : n10534_o;
  assign n10536_o = n9735_o[1007:1000];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10537_o = n10155_o ? wdata_i : n10536_o;
  assign n10538_o = n9735_o[1015:1008];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10539_o = n10156_o ? wdata_i : n10538_o;
  assign n10540_o = n9735_o[1023:1016];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10541_o = n10157_o ? wdata_i : n10540_o;
  assign n10542_o = n9735_o[1031:1024];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10543_o = n10158_o ? wdata_i : n10542_o;
  assign n10544_o = n9735_o[1039:1032];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10545_o = n10159_o ? wdata_i : n10544_o;
  assign n10546_o = n9735_o[1047:1040];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10547_o = n10160_o ? wdata_i : n10546_o;
  assign n10548_o = n9735_o[1055:1048];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10549_o = n10161_o ? wdata_i : n10548_o;
  assign n10550_o = n9735_o[1063:1056];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10551_o = n10162_o ? wdata_i : n10550_o;
  assign n10552_o = n9735_o[1071:1064];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10553_o = n10163_o ? wdata_i : n10552_o;
  assign n10554_o = n9735_o[1079:1072];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10555_o = n10164_o ? wdata_i : n10554_o;
  assign n10556_o = n9735_o[1087:1080];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10557_o = n10165_o ? wdata_i : n10556_o;
  assign n10558_o = n9735_o[1095:1088];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10559_o = n10166_o ? wdata_i : n10558_o;
  assign n10560_o = n9735_o[1103:1096];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10561_o = n10167_o ? wdata_i : n10560_o;
  assign n10562_o = n9735_o[1111:1104];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10563_o = n10168_o ? wdata_i : n10562_o;
  assign n10564_o = n9735_o[1119:1112];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10565_o = n10169_o ? wdata_i : n10564_o;
  assign n10566_o = n9735_o[1127:1120];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10567_o = n10170_o ? wdata_i : n10566_o;
  assign n10568_o = n9735_o[1135:1128];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10569_o = n10171_o ? wdata_i : n10568_o;
  assign n10570_o = n9735_o[1143:1136];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10571_o = n10172_o ? wdata_i : n10570_o;
  assign n10572_o = n9735_o[1151:1144];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10573_o = n10173_o ? wdata_i : n10572_o;
  assign n10574_o = n9735_o[1159:1152];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10575_o = n10174_o ? wdata_i : n10574_o;
  assign n10576_o = n9735_o[1167:1160];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10577_o = n10175_o ? wdata_i : n10576_o;
  assign n10578_o = n9735_o[1175:1168];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10579_o = n10176_o ? wdata_i : n10578_o;
  assign n10580_o = n9735_o[1183:1176];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10581_o = n10177_o ? wdata_i : n10580_o;
  assign n10582_o = n9735_o[1191:1184];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10583_o = n10178_o ? wdata_i : n10582_o;
  assign n10584_o = n9735_o[1199:1192];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10585_o = n10179_o ? wdata_i : n10584_o;
  assign n10586_o = n9735_o[1207:1200];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10587_o = n10180_o ? wdata_i : n10586_o;
  assign n10588_o = n9735_o[1215:1208];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10589_o = n10181_o ? wdata_i : n10588_o;
  assign n10590_o = n9735_o[1223:1216];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10591_o = n10182_o ? wdata_i : n10590_o;
  assign n10592_o = n9735_o[1231:1224];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10593_o = n10183_o ? wdata_i : n10592_o;
  assign n10594_o = n9735_o[1239:1232];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10595_o = n10184_o ? wdata_i : n10594_o;
  assign n10596_o = n9735_o[1247:1240];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10597_o = n10185_o ? wdata_i : n10596_o;
  assign n10598_o = n9735_o[1255:1248];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10599_o = n10186_o ? wdata_i : n10598_o;
  assign n10600_o = n9735_o[1263:1256];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10601_o = n10187_o ? wdata_i : n10600_o;
  assign n10602_o = n9735_o[1271:1264];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10603_o = n10188_o ? wdata_i : n10602_o;
  assign n10604_o = n9735_o[1279:1272];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10605_o = n10189_o ? wdata_i : n10604_o;
  assign n10606_o = n9735_o[1287:1280];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10607_o = n10190_o ? wdata_i : n10606_o;
  assign n10608_o = n9735_o[1295:1288];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10609_o = n10191_o ? wdata_i : n10608_o;
  assign n10610_o = n9735_o[1303:1296];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10611_o = n10192_o ? wdata_i : n10610_o;
  assign n10612_o = n9735_o[1311:1304];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10613_o = n10193_o ? wdata_i : n10612_o;
  assign n10614_o = n9735_o[1319:1312];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10615_o = n10194_o ? wdata_i : n10614_o;
  assign n10616_o = n9735_o[1327:1320];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10617_o = n10195_o ? wdata_i : n10616_o;
  assign n10618_o = n9735_o[1335:1328];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10619_o = n10196_o ? wdata_i : n10618_o;
  assign n10620_o = n9735_o[1343:1336];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10621_o = n10197_o ? wdata_i : n10620_o;
  assign n10622_o = n9735_o[1351:1344];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10623_o = n10198_o ? wdata_i : n10622_o;
  assign n10624_o = n9735_o[1359:1352];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10625_o = n10199_o ? wdata_i : n10624_o;
  assign n10626_o = n9735_o[1367:1360];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10627_o = n10200_o ? wdata_i : n10626_o;
  assign n10628_o = n9735_o[1375:1368];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10629_o = n10201_o ? wdata_i : n10628_o;
  assign n10630_o = n9735_o[1383:1376];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10631_o = n10202_o ? wdata_i : n10630_o;
  assign n10632_o = n9735_o[1391:1384];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10633_o = n10203_o ? wdata_i : n10632_o;
  assign n10634_o = n9735_o[1399:1392];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10635_o = n10204_o ? wdata_i : n10634_o;
  assign n10636_o = n9735_o[1407:1400];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10637_o = n10205_o ? wdata_i : n10636_o;
  assign n10638_o = n9735_o[1415:1408];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10639_o = n10206_o ? wdata_i : n10638_o;
  assign n10640_o = n9735_o[1423:1416];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10641_o = n10207_o ? wdata_i : n10640_o;
  assign n10642_o = n9735_o[1431:1424];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10643_o = n10208_o ? wdata_i : n10642_o;
  assign n10644_o = n9735_o[1439:1432];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10645_o = n10209_o ? wdata_i : n10644_o;
  assign n10646_o = n9735_o[1447:1440];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10647_o = n10210_o ? wdata_i : n10646_o;
  assign n10648_o = n9735_o[1455:1448];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10649_o = n10211_o ? wdata_i : n10648_o;
  assign n10650_o = n9735_o[1463:1456];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10651_o = n10212_o ? wdata_i : n10650_o;
  assign n10652_o = n9735_o[1471:1464];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10653_o = n10213_o ? wdata_i : n10652_o;
  assign n10654_o = n9735_o[1479:1472];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10655_o = n10214_o ? wdata_i : n10654_o;
  assign n10656_o = n9735_o[1487:1480];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10657_o = n10215_o ? wdata_i : n10656_o;
  assign n10658_o = n9735_o[1495:1488];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10659_o = n10216_o ? wdata_i : n10658_o;
  assign n10660_o = n9735_o[1503:1496];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10661_o = n10217_o ? wdata_i : n10660_o;
  assign n10662_o = n9735_o[1511:1504];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10663_o = n10218_o ? wdata_i : n10662_o;
  assign n10664_o = n9735_o[1519:1512];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10665_o = n10219_o ? wdata_i : n10664_o;
  assign n10666_o = n9735_o[1527:1520];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10667_o = n10220_o ? wdata_i : n10666_o;
  assign n10668_o = n9735_o[1535:1528];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10669_o = n10221_o ? wdata_i : n10668_o;
  assign n10670_o = n9735_o[1543:1536];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10671_o = n10222_o ? wdata_i : n10670_o;
  assign n10672_o = n9735_o[1551:1544];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10673_o = n10223_o ? wdata_i : n10672_o;
  assign n10674_o = n9735_o[1559:1552];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10675_o = n10224_o ? wdata_i : n10674_o;
  assign n10676_o = n9735_o[1567:1560];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10677_o = n10225_o ? wdata_i : n10676_o;
  assign n10678_o = n9735_o[1575:1568];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10679_o = n10226_o ? wdata_i : n10678_o;
  assign n10680_o = n9735_o[1583:1576];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10681_o = n10227_o ? wdata_i : n10680_o;
  assign n10682_o = n9735_o[1591:1584];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10683_o = n10228_o ? wdata_i : n10682_o;
  assign n10684_o = n9735_o[1599:1592];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10685_o = n10229_o ? wdata_i : n10684_o;
  assign n10686_o = n9735_o[1607:1600];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10687_o = n10230_o ? wdata_i : n10686_o;
  assign n10688_o = n9735_o[1615:1608];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10689_o = n10231_o ? wdata_i : n10688_o;
  assign n10690_o = n9735_o[1623:1616];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10691_o = n10232_o ? wdata_i : n10690_o;
  assign n10692_o = n9735_o[1631:1624];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10693_o = n10233_o ? wdata_i : n10692_o;
  assign n10694_o = n9735_o[1639:1632];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10695_o = n10234_o ? wdata_i : n10694_o;
  assign n10696_o = n9735_o[1647:1640];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10697_o = n10235_o ? wdata_i : n10696_o;
  assign n10698_o = n9735_o[1655:1648];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10699_o = n10236_o ? wdata_i : n10698_o;
  assign n10700_o = n9735_o[1663:1656];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10701_o = n10237_o ? wdata_i : n10700_o;
  assign n10702_o = n9735_o[1671:1664];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10703_o = n10238_o ? wdata_i : n10702_o;
  assign n10704_o = n9735_o[1679:1672];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10705_o = n10239_o ? wdata_i : n10704_o;
  assign n10706_o = n9735_o[1687:1680];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10707_o = n10240_o ? wdata_i : n10706_o;
  assign n10708_o = n9735_o[1695:1688];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10709_o = n10241_o ? wdata_i : n10708_o;
  assign n10710_o = n9735_o[1703:1696];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10711_o = n10242_o ? wdata_i : n10710_o;
  assign n10712_o = n9735_o[1711:1704];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10713_o = n10243_o ? wdata_i : n10712_o;
  assign n10714_o = n9735_o[1719:1712];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10715_o = n10244_o ? wdata_i : n10714_o;
  assign n10716_o = n9735_o[1727:1720];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10717_o = n10245_o ? wdata_i : n10716_o;
  assign n10718_o = n9735_o[1735:1728];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10719_o = n10246_o ? wdata_i : n10718_o;
  assign n10720_o = n9735_o[1743:1736];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10721_o = n10247_o ? wdata_i : n10720_o;
  assign n10722_o = n9735_o[1751:1744];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10723_o = n10248_o ? wdata_i : n10722_o;
  assign n10724_o = n9735_o[1759:1752];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10725_o = n10249_o ? wdata_i : n10724_o;
  assign n10726_o = n9735_o[1767:1760];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10727_o = n10250_o ? wdata_i : n10726_o;
  assign n10728_o = n9735_o[1775:1768];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10729_o = n10251_o ? wdata_i : n10728_o;
  assign n10730_o = n9735_o[1783:1776];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10731_o = n10252_o ? wdata_i : n10730_o;
  assign n10732_o = n9735_o[1791:1784];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10733_o = n10253_o ? wdata_i : n10732_o;
  assign n10734_o = n9735_o[1799:1792];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10735_o = n10254_o ? wdata_i : n10734_o;
  assign n10736_o = n9735_o[1807:1800];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10737_o = n10255_o ? wdata_i : n10736_o;
  assign n10738_o = n9735_o[1815:1808];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10739_o = n10256_o ? wdata_i : n10738_o;
  assign n10740_o = n9735_o[1823:1816];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10741_o = n10257_o ? wdata_i : n10740_o;
  assign n10742_o = n9735_o[1831:1824];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10743_o = n10258_o ? wdata_i : n10742_o;
  assign n10744_o = n9735_o[1839:1832];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10745_o = n10259_o ? wdata_i : n10744_o;
  assign n10746_o = n9735_o[1847:1840];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10747_o = n10260_o ? wdata_i : n10746_o;
  assign n10748_o = n9735_o[1855:1848];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10749_o = n10261_o ? wdata_i : n10748_o;
  assign n10750_o = n9735_o[1863:1856];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10751_o = n10262_o ? wdata_i : n10750_o;
  assign n10752_o = n9735_o[1871:1864];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10753_o = n10263_o ? wdata_i : n10752_o;
  assign n10754_o = n9735_o[1879:1872];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10755_o = n10264_o ? wdata_i : n10754_o;
  assign n10756_o = n9735_o[1887:1880];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10757_o = n10265_o ? wdata_i : n10756_o;
  assign n10758_o = n9735_o[1895:1888];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10759_o = n10266_o ? wdata_i : n10758_o;
  assign n10760_o = n9735_o[1903:1896];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10761_o = n10267_o ? wdata_i : n10760_o;
  assign n10762_o = n9735_o[1911:1904];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10763_o = n10268_o ? wdata_i : n10762_o;
  assign n10764_o = n9735_o[1919:1912];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10765_o = n10269_o ? wdata_i : n10764_o;
  assign n10766_o = n9735_o[1927:1920];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10767_o = n10270_o ? wdata_i : n10766_o;
  assign n10768_o = n9735_o[1935:1928];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10769_o = n10271_o ? wdata_i : n10768_o;
  assign n10770_o = n9735_o[1943:1936];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10771_o = n10272_o ? wdata_i : n10770_o;
  assign n10772_o = n9735_o[1951:1944];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10773_o = n10273_o ? wdata_i : n10772_o;
  assign n10774_o = n9735_o[1959:1952];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10775_o = n10274_o ? wdata_i : n10774_o;
  assign n10776_o = n9735_o[1967:1960];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10777_o = n10275_o ? wdata_i : n10776_o;
  assign n10778_o = n9735_o[1975:1968];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10779_o = n10276_o ? wdata_i : n10778_o;
  assign n10780_o = n9735_o[1983:1976];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10781_o = n10277_o ? wdata_i : n10780_o;
  assign n10782_o = n9735_o[1991:1984];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10783_o = n10278_o ? wdata_i : n10782_o;
  assign n10784_o = n9735_o[1999:1992];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10785_o = n10279_o ? wdata_i : n10784_o;
  assign n10786_o = n9735_o[2007:2000];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10787_o = n10280_o ? wdata_i : n10786_o;
  assign n10788_o = n9735_o[2015:2008];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10789_o = n10281_o ? wdata_i : n10788_o;
  assign n10790_o = n9735_o[2023:2016];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10791_o = n10282_o ? wdata_i : n10790_o;
  assign n10792_o = n9735_o[2031:2024];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10793_o = n10283_o ? wdata_i : n10792_o;
  assign n10794_o = n9735_o[2039:2032];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10795_o = n10284_o ? wdata_i : n10794_o;
  assign n10796_o = n9735_o[2047:2040];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10797_o = n10285_o ? wdata_i : n10796_o;
  assign n10798_o = {n10797_o, n10795_o, n10793_o, n10791_o, n10789_o, n10787_o, n10785_o, n10783_o, n10781_o, n10779_o, n10777_o, n10775_o, n10773_o, n10771_o, n10769_o, n10767_o, n10765_o, n10763_o, n10761_o, n10759_o, n10757_o, n10755_o, n10753_o, n10751_o, n10749_o, n10747_o, n10745_o, n10743_o, n10741_o, n10739_o, n10737_o, n10735_o, n10733_o, n10731_o, n10729_o, n10727_o, n10725_o, n10723_o, n10721_o, n10719_o, n10717_o, n10715_o, n10713_o, n10711_o, n10709_o, n10707_o, n10705_o, n10703_o, n10701_o, n10699_o, n10697_o, n10695_o, n10693_o, n10691_o, n10689_o, n10687_o, n10685_o, n10683_o, n10681_o, n10679_o, n10677_o, n10675_o, n10673_o, n10671_o, n10669_o, n10667_o, n10665_o, n10663_o, n10661_o, n10659_o, n10657_o, n10655_o, n10653_o, n10651_o, n10649_o, n10647_o, n10645_o, n10643_o, n10641_o, n10639_o, n10637_o, n10635_o, n10633_o, n10631_o, n10629_o, n10627_o, n10625_o, n10623_o, n10621_o, n10619_o, n10617_o, n10615_o, n10613_o, n10611_o, n10609_o, n10607_o, n10605_o, n10603_o, n10601_o, n10599_o, n10597_o, n10595_o, n10593_o, n10591_o, n10589_o, n10587_o, n10585_o, n10583_o, n10581_o, n10579_o, n10577_o, n10575_o, n10573_o, n10571_o, n10569_o, n10567_o, n10565_o, n10563_o, n10561_o, n10559_o, n10557_o, n10555_o, n10553_o, n10551_o, n10549_o, n10547_o, n10545_o, n10543_o, n10541_o, n10539_o, n10537_o, n10535_o, n10533_o, n10531_o, n10529_o, n10527_o, n10525_o, n10523_o, n10521_o, n10519_o, n10517_o, n10515_o, n10513_o, n10511_o, n10509_o, n10507_o, n10505_o, n10503_o, n10501_o, n10499_o, n10497_o, n10495_o, n10493_o, n10491_o, n10489_o, n10487_o, n10485_o, n10483_o, n10481_o, n10479_o, n10477_o, n10475_o, n10473_o, n10471_o, n10469_o, n10467_o, n10465_o, n10463_o, n10461_o, n10459_o, n10457_o, n10455_o, n10453_o, n10451_o, n10449_o, n10447_o, n10445_o, n10443_o, n10441_o, n10439_o, n10437_o, n10435_o, n10433_o, n10431_o, n10429_o, n10427_o, n10425_o, n10423_o, n10421_o, n10419_o, n10417_o, n10415_o, n10413_o, n10411_o, n10409_o, n10407_o, n10405_o, n10403_o, n10401_o, n10399_o, n10397_o, n10395_o, n10393_o, n10391_o, n10389_o, n10387_o, n10385_o, n10383_o, n10381_o, n10379_o, n10377_o, n10375_o, n10373_o, n10371_o, n10369_o, n10367_o, n10365_o, n10363_o, n10361_o, n10359_o, n10357_o, n10355_o, n10353_o, n10351_o, n10349_o, n10347_o, n10345_o, n10343_o, n10341_o, n10339_o, n10337_o, n10335_o, n10333_o, n10331_o, n10329_o, n10327_o, n10325_o, n10323_o, n10321_o, n10319_o, n10317_o, n10315_o, n10313_o, n10311_o, n10309_o, n10307_o, n10305_o, n10303_o, n10301_o, n10299_o, n10297_o, n10295_o, n10293_o, n10291_o, n10289_o, n10287_o};
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:21  */
  assign n10799_o = fifo[27:20];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:184:11  */
  assign n10800_o = fifo[35:28];
  assign n10801_o = fifo[43:36];
  assign n10802_o = fifo[51:44];
  assign n10803_o = fifo[59:52];
  assign n10804_o = fifo[67:60];
  assign n10805_o = fifo[75:68];
  assign n10806_o = fifo[83:76];
  assign n10807_o = fifo[91:84];
  assign n10808_o = fifo[99:92];
  assign n10809_o = fifo[107:100];
  assign n10810_o = fifo[115:108];
  assign n10811_o = fifo[123:116];
  assign n10812_o = fifo[131:124];
  assign n10813_o = fifo[139:132];
  assign n10814_o = fifo[147:140];
  assign n10815_o = fifo[155:148];
  assign n10816_o = fifo[163:156];
  assign n10817_o = fifo[171:164];
  assign n10818_o = fifo[179:172];
  assign n10819_o = fifo[187:180];
  assign n10820_o = fifo[195:188];
  assign n10821_o = fifo[203:196];
  assign n10822_o = fifo[211:204];
  assign n10823_o = fifo[219:212];
  assign n10824_o = fifo[227:220];
  assign n10825_o = fifo[235:228];
  assign n10826_o = fifo[243:236];
  assign n10827_o = fifo[251:244];
  assign n10828_o = fifo[259:252];
  assign n10829_o = fifo[267:260];
  assign n10830_o = fifo[275:268];
  assign n10831_o = fifo[283:276];
  assign n10832_o = fifo[291:284];
  assign n10833_o = fifo[299:292];
  assign n10834_o = fifo[307:300];
  assign n10835_o = fifo[315:308];
  assign n10836_o = fifo[323:316];
  assign n10837_o = fifo[331:324];
  assign n10838_o = fifo[339:332];
  assign n10839_o = fifo[347:340];
  assign n10840_o = fifo[355:348];
  assign n10841_o = fifo[363:356];
  assign n10842_o = fifo[371:364];
  assign n10843_o = fifo[379:372];
  assign n10844_o = fifo[387:380];
  assign n10845_o = fifo[395:388];
  assign n10846_o = fifo[403:396];
  assign n10847_o = fifo[411:404];
  assign n10848_o = fifo[419:412];
  assign n10849_o = fifo[427:420];
  assign n10850_o = fifo[435:428];
  assign n10851_o = fifo[443:436];
  assign n10852_o = fifo[451:444];
  assign n10853_o = fifo[459:452];
  assign n10854_o = fifo[467:460];
  assign n10855_o = fifo[475:468];
  assign n10856_o = fifo[483:476];
  assign n10857_o = fifo[491:484];
  assign n10858_o = fifo[499:492];
  assign n10859_o = fifo[507:500];
  assign n10860_o = fifo[515:508];
  assign n10861_o = fifo[523:516];
  assign n10862_o = fifo[531:524];
  assign n10863_o = fifo[539:532];
  assign n10864_o = fifo[547:540];
  assign n10865_o = fifo[555:548];
  assign n10866_o = fifo[563:556];
  assign n10867_o = fifo[571:564];
  assign n10868_o = fifo[579:572];
  assign n10869_o = fifo[587:580];
  assign n10870_o = fifo[595:588];
  assign n10871_o = fifo[603:596];
  assign n10872_o = fifo[611:604];
  assign n10873_o = fifo[619:612];
  assign n10874_o = fifo[627:620];
  assign n10875_o = fifo[635:628];
  assign n10876_o = fifo[643:636];
  assign n10877_o = fifo[651:644];
  assign n10878_o = fifo[659:652];
  assign n10879_o = fifo[667:660];
  assign n10880_o = fifo[675:668];
  assign n10881_o = fifo[683:676];
  assign n10882_o = fifo[691:684];
  assign n10883_o = fifo[699:692];
  assign n10884_o = fifo[707:700];
  assign n10885_o = fifo[715:708];
  assign n10886_o = fifo[723:716];
  assign n10887_o = fifo[731:724];
  assign n10888_o = fifo[739:732];
  assign n10889_o = fifo[747:740];
  assign n10890_o = fifo[755:748];
  assign n10891_o = fifo[763:756];
  assign n10892_o = fifo[771:764];
  assign n10893_o = fifo[779:772];
  assign n10894_o = fifo[787:780];
  assign n10895_o = fifo[795:788];
  assign n10896_o = fifo[803:796];
  assign n10897_o = fifo[811:804];
  assign n10898_o = fifo[819:812];
  assign n10899_o = fifo[827:820];
  assign n10900_o = fifo[835:828];
  assign n10901_o = fifo[843:836];
  assign n10902_o = fifo[851:844];
  assign n10903_o = fifo[859:852];
  assign n10904_o = fifo[867:860];
  assign n10905_o = fifo[875:868];
  assign n10906_o = fifo[883:876];
  assign n10907_o = fifo[891:884];
  assign n10908_o = fifo[899:892];
  assign n10909_o = fifo[907:900];
  assign n10910_o = fifo[915:908];
  assign n10911_o = fifo[923:916];
  assign n10912_o = fifo[931:924];
  assign n10913_o = fifo[939:932];
  assign n10914_o = fifo[947:940];
  assign n10915_o = fifo[955:948];
  assign n10916_o = fifo[963:956];
  assign n10917_o = fifo[971:964];
  assign n10918_o = fifo[979:972];
  assign n10919_o = fifo[987:980];
  assign n10920_o = fifo[995:988];
  assign n10921_o = fifo[1003:996];
  assign n10922_o = fifo[1011:1004];
  assign n10923_o = fifo[1019:1012];
  assign n10924_o = fifo[1027:1020];
  assign n10925_o = fifo[1035:1028];
  assign n10926_o = fifo[1043:1036];
  assign n10927_o = fifo[1051:1044];
  assign n10928_o = fifo[1059:1052];
  assign n10929_o = fifo[1067:1060];
  assign n10930_o = fifo[1075:1068];
  assign n10931_o = fifo[1083:1076];
  assign n10932_o = fifo[1091:1084];
  assign n10933_o = fifo[1099:1092];
  assign n10934_o = fifo[1107:1100];
  assign n10935_o = fifo[1115:1108];
  assign n10936_o = fifo[1123:1116];
  assign n10937_o = fifo[1131:1124];
  assign n10938_o = fifo[1139:1132];
  assign n10939_o = fifo[1147:1140];
  assign n10940_o = fifo[1155:1148];
  assign n10941_o = fifo[1163:1156];
  assign n10942_o = fifo[1171:1164];
  assign n10943_o = fifo[1179:1172];
  assign n10944_o = fifo[1187:1180];
  assign n10945_o = fifo[1195:1188];
  assign n10946_o = fifo[1203:1196];
  assign n10947_o = fifo[1211:1204];
  assign n10948_o = fifo[1219:1212];
  assign n10949_o = fifo[1227:1220];
  assign n10950_o = fifo[1235:1228];
  assign n10951_o = fifo[1243:1236];
  assign n10952_o = fifo[1251:1244];
  assign n10953_o = fifo[1259:1252];
  assign n10954_o = fifo[1267:1260];
  assign n10955_o = fifo[1275:1268];
  assign n10956_o = fifo[1283:1276];
  assign n10957_o = fifo[1291:1284];
  assign n10958_o = fifo[1299:1292];
  assign n10959_o = fifo[1307:1300];
  assign n10960_o = fifo[1315:1308];
  assign n10961_o = fifo[1323:1316];
  assign n10962_o = fifo[1331:1324];
  assign n10963_o = fifo[1339:1332];
  assign n10964_o = fifo[1347:1340];
  assign n10965_o = fifo[1355:1348];
  assign n10966_o = fifo[1363:1356];
  assign n10967_o = fifo[1371:1364];
  assign n10968_o = fifo[1379:1372];
  assign n10969_o = fifo[1387:1380];
  assign n10970_o = fifo[1395:1388];
  assign n10971_o = fifo[1403:1396];
  assign n10972_o = fifo[1411:1404];
  assign n10973_o = fifo[1419:1412];
  assign n10974_o = fifo[1427:1420];
  assign n10975_o = fifo[1435:1428];
  assign n10976_o = fifo[1443:1436];
  assign n10977_o = fifo[1451:1444];
  assign n10978_o = fifo[1459:1452];
  assign n10979_o = fifo[1467:1460];
  assign n10980_o = fifo[1475:1468];
  assign n10981_o = fifo[1483:1476];
  assign n10982_o = fifo[1491:1484];
  assign n10983_o = fifo[1499:1492];
  assign n10984_o = fifo[1507:1500];
  assign n10985_o = fifo[1515:1508];
  assign n10986_o = fifo[1523:1516];
  assign n10987_o = fifo[1531:1524];
  assign n10988_o = fifo[1539:1532];
  assign n10989_o = fifo[1547:1540];
  assign n10990_o = fifo[1555:1548];
  assign n10991_o = fifo[1563:1556];
  assign n10992_o = fifo[1571:1564];
  assign n10993_o = fifo[1579:1572];
  assign n10994_o = fifo[1587:1580];
  assign n10995_o = fifo[1595:1588];
  assign n10996_o = fifo[1603:1596];
  assign n10997_o = fifo[1611:1604];
  assign n10998_o = fifo[1619:1612];
  assign n10999_o = fifo[1627:1620];
  assign n11000_o = fifo[1635:1628];
  assign n11001_o = fifo[1643:1636];
  assign n11002_o = fifo[1651:1644];
  assign n11003_o = fifo[1659:1652];
  assign n11004_o = fifo[1667:1660];
  assign n11005_o = fifo[1675:1668];
  assign n11006_o = fifo[1683:1676];
  assign n11007_o = fifo[1691:1684];
  assign n11008_o = fifo[1699:1692];
  assign n11009_o = fifo[1707:1700];
  assign n11010_o = fifo[1715:1708];
  assign n11011_o = fifo[1723:1716];
  assign n11012_o = fifo[1731:1724];
  assign n11013_o = fifo[1739:1732];
  assign n11014_o = fifo[1747:1740];
  assign n11015_o = fifo[1755:1748];
  assign n11016_o = fifo[1763:1756];
  assign n11017_o = fifo[1771:1764];
  assign n11018_o = fifo[1779:1772];
  assign n11019_o = fifo[1787:1780];
  assign n11020_o = fifo[1795:1788];
  assign n11021_o = fifo[1803:1796];
  assign n11022_o = fifo[1811:1804];
  assign n11023_o = fifo[1819:1812];
  assign n11024_o = fifo[1827:1820];
  assign n11025_o = fifo[1835:1828];
  assign n11026_o = fifo[1843:1836];
  assign n11027_o = fifo[1851:1844];
  assign n11028_o = fifo[1859:1852];
  assign n11029_o = fifo[1867:1860];
  assign n11030_o = fifo[1875:1868];
  assign n11031_o = fifo[1883:1876];
  assign n11032_o = fifo[1891:1884];
  assign n11033_o = fifo[1899:1892];
  assign n11034_o = fifo[1907:1900];
  assign n11035_o = fifo[1915:1908];
  assign n11036_o = fifo[1923:1916];
  assign n11037_o = fifo[1931:1924];
  assign n11038_o = fifo[1939:1932];
  assign n11039_o = fifo[1947:1940];
  assign n11040_o = fifo[1955:1948];
  assign n11041_o = fifo[1963:1956];
  assign n11042_o = fifo[1971:1964];
  assign n11043_o = fifo[1979:1972];
  assign n11044_o = fifo[1987:1980];
  assign n11045_o = fifo[1995:1988];
  assign n11046_o = fifo[2003:1996];
  assign n11047_o = fifo[2011:2004];
  assign n11048_o = fifo[2019:2012];
  assign n11049_o = fifo[2027:2020];
  assign n11050_o = fifo[2035:2028];
  assign n11051_o = fifo[2043:2036];
  assign n11052_o = fifo[2051:2044];
  assign n11053_o = fifo[2059:2052];
  assign n11054_o = fifo[2067:2060];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11055_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11055_o)
      2'b00: n11056_o = n10799_o;
      2'b01: n11056_o = n10800_o;
      2'b10: n11056_o = n10801_o;
      2'b11: n11056_o = n10802_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11057_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11057_o)
      2'b00: n11058_o = n10803_o;
      2'b01: n11058_o = n10804_o;
      2'b10: n11058_o = n10805_o;
      2'b11: n11058_o = n10806_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11059_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11059_o)
      2'b00: n11060_o = n10807_o;
      2'b01: n11060_o = n10808_o;
      2'b10: n11060_o = n10809_o;
      2'b11: n11060_o = n10810_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11061_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11061_o)
      2'b00: n11062_o = n10811_o;
      2'b01: n11062_o = n10812_o;
      2'b10: n11062_o = n10813_o;
      2'b11: n11062_o = n10814_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11063_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11063_o)
      2'b00: n11064_o = n10815_o;
      2'b01: n11064_o = n10816_o;
      2'b10: n11064_o = n10817_o;
      2'b11: n11064_o = n10818_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11065_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11065_o)
      2'b00: n11066_o = n10819_o;
      2'b01: n11066_o = n10820_o;
      2'b10: n11066_o = n10821_o;
      2'b11: n11066_o = n10822_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11067_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11067_o)
      2'b00: n11068_o = n10823_o;
      2'b01: n11068_o = n10824_o;
      2'b10: n11068_o = n10825_o;
      2'b11: n11068_o = n10826_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11069_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11069_o)
      2'b00: n11070_o = n10827_o;
      2'b01: n11070_o = n10828_o;
      2'b10: n11070_o = n10829_o;
      2'b11: n11070_o = n10830_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11071_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11071_o)
      2'b00: n11072_o = n10831_o;
      2'b01: n11072_o = n10832_o;
      2'b10: n11072_o = n10833_o;
      2'b11: n11072_o = n10834_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11073_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11073_o)
      2'b00: n11074_o = n10835_o;
      2'b01: n11074_o = n10836_o;
      2'b10: n11074_o = n10837_o;
      2'b11: n11074_o = n10838_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11075_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11075_o)
      2'b00: n11076_o = n10839_o;
      2'b01: n11076_o = n10840_o;
      2'b10: n11076_o = n10841_o;
      2'b11: n11076_o = n10842_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11077_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11077_o)
      2'b00: n11078_o = n10843_o;
      2'b01: n11078_o = n10844_o;
      2'b10: n11078_o = n10845_o;
      2'b11: n11078_o = n10846_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11079_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11079_o)
      2'b00: n11080_o = n10847_o;
      2'b01: n11080_o = n10848_o;
      2'b10: n11080_o = n10849_o;
      2'b11: n11080_o = n10850_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11081_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11081_o)
      2'b00: n11082_o = n10851_o;
      2'b01: n11082_o = n10852_o;
      2'b10: n11082_o = n10853_o;
      2'b11: n11082_o = n10854_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11083_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11083_o)
      2'b00: n11084_o = n10855_o;
      2'b01: n11084_o = n10856_o;
      2'b10: n11084_o = n10857_o;
      2'b11: n11084_o = n10858_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11085_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11085_o)
      2'b00: n11086_o = n10859_o;
      2'b01: n11086_o = n10860_o;
      2'b10: n11086_o = n10861_o;
      2'b11: n11086_o = n10862_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11087_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11087_o)
      2'b00: n11088_o = n10863_o;
      2'b01: n11088_o = n10864_o;
      2'b10: n11088_o = n10865_o;
      2'b11: n11088_o = n10866_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11089_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11089_o)
      2'b00: n11090_o = n10867_o;
      2'b01: n11090_o = n10868_o;
      2'b10: n11090_o = n10869_o;
      2'b11: n11090_o = n10870_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11091_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11091_o)
      2'b00: n11092_o = n10871_o;
      2'b01: n11092_o = n10872_o;
      2'b10: n11092_o = n10873_o;
      2'b11: n11092_o = n10874_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11093_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11093_o)
      2'b00: n11094_o = n10875_o;
      2'b01: n11094_o = n10876_o;
      2'b10: n11094_o = n10877_o;
      2'b11: n11094_o = n10878_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11095_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11095_o)
      2'b00: n11096_o = n10879_o;
      2'b01: n11096_o = n10880_o;
      2'b10: n11096_o = n10881_o;
      2'b11: n11096_o = n10882_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11097_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11097_o)
      2'b00: n11098_o = n10883_o;
      2'b01: n11098_o = n10884_o;
      2'b10: n11098_o = n10885_o;
      2'b11: n11098_o = n10886_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11099_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11099_o)
      2'b00: n11100_o = n10887_o;
      2'b01: n11100_o = n10888_o;
      2'b10: n11100_o = n10889_o;
      2'b11: n11100_o = n10890_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11101_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11101_o)
      2'b00: n11102_o = n10891_o;
      2'b01: n11102_o = n10892_o;
      2'b10: n11102_o = n10893_o;
      2'b11: n11102_o = n10894_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11103_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11103_o)
      2'b00: n11104_o = n10895_o;
      2'b01: n11104_o = n10896_o;
      2'b10: n11104_o = n10897_o;
      2'b11: n11104_o = n10898_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11105_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11105_o)
      2'b00: n11106_o = n10899_o;
      2'b01: n11106_o = n10900_o;
      2'b10: n11106_o = n10901_o;
      2'b11: n11106_o = n10902_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11107_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11107_o)
      2'b00: n11108_o = n10903_o;
      2'b01: n11108_o = n10904_o;
      2'b10: n11108_o = n10905_o;
      2'b11: n11108_o = n10906_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11109_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11109_o)
      2'b00: n11110_o = n10907_o;
      2'b01: n11110_o = n10908_o;
      2'b10: n11110_o = n10909_o;
      2'b11: n11110_o = n10910_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11111_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11111_o)
      2'b00: n11112_o = n10911_o;
      2'b01: n11112_o = n10912_o;
      2'b10: n11112_o = n10913_o;
      2'b11: n11112_o = n10914_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11113_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11113_o)
      2'b00: n11114_o = n10915_o;
      2'b01: n11114_o = n10916_o;
      2'b10: n11114_o = n10917_o;
      2'b11: n11114_o = n10918_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11115_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11115_o)
      2'b00: n11116_o = n10919_o;
      2'b01: n11116_o = n10920_o;
      2'b10: n11116_o = n10921_o;
      2'b11: n11116_o = n10922_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11117_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11117_o)
      2'b00: n11118_o = n10923_o;
      2'b01: n11118_o = n10924_o;
      2'b10: n11118_o = n10925_o;
      2'b11: n11118_o = n10926_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11119_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11119_o)
      2'b00: n11120_o = n10927_o;
      2'b01: n11120_o = n10928_o;
      2'b10: n11120_o = n10929_o;
      2'b11: n11120_o = n10930_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11121_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11121_o)
      2'b00: n11122_o = n10931_o;
      2'b01: n11122_o = n10932_o;
      2'b10: n11122_o = n10933_o;
      2'b11: n11122_o = n10934_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11123_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11123_o)
      2'b00: n11124_o = n10935_o;
      2'b01: n11124_o = n10936_o;
      2'b10: n11124_o = n10937_o;
      2'b11: n11124_o = n10938_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11125_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11125_o)
      2'b00: n11126_o = n10939_o;
      2'b01: n11126_o = n10940_o;
      2'b10: n11126_o = n10941_o;
      2'b11: n11126_o = n10942_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11127_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11127_o)
      2'b00: n11128_o = n10943_o;
      2'b01: n11128_o = n10944_o;
      2'b10: n11128_o = n10945_o;
      2'b11: n11128_o = n10946_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11129_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11129_o)
      2'b00: n11130_o = n10947_o;
      2'b01: n11130_o = n10948_o;
      2'b10: n11130_o = n10949_o;
      2'b11: n11130_o = n10950_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11131_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11131_o)
      2'b00: n11132_o = n10951_o;
      2'b01: n11132_o = n10952_o;
      2'b10: n11132_o = n10953_o;
      2'b11: n11132_o = n10954_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11133_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11133_o)
      2'b00: n11134_o = n10955_o;
      2'b01: n11134_o = n10956_o;
      2'b10: n11134_o = n10957_o;
      2'b11: n11134_o = n10958_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11135_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11135_o)
      2'b00: n11136_o = n10959_o;
      2'b01: n11136_o = n10960_o;
      2'b10: n11136_o = n10961_o;
      2'b11: n11136_o = n10962_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11137_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11137_o)
      2'b00: n11138_o = n10963_o;
      2'b01: n11138_o = n10964_o;
      2'b10: n11138_o = n10965_o;
      2'b11: n11138_o = n10966_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11139_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11139_o)
      2'b00: n11140_o = n10967_o;
      2'b01: n11140_o = n10968_o;
      2'b10: n11140_o = n10969_o;
      2'b11: n11140_o = n10970_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11141_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11141_o)
      2'b00: n11142_o = n10971_o;
      2'b01: n11142_o = n10972_o;
      2'b10: n11142_o = n10973_o;
      2'b11: n11142_o = n10974_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11143_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11143_o)
      2'b00: n11144_o = n10975_o;
      2'b01: n11144_o = n10976_o;
      2'b10: n11144_o = n10977_o;
      2'b11: n11144_o = n10978_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11145_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11145_o)
      2'b00: n11146_o = n10979_o;
      2'b01: n11146_o = n10980_o;
      2'b10: n11146_o = n10981_o;
      2'b11: n11146_o = n10982_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11147_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11147_o)
      2'b00: n11148_o = n10983_o;
      2'b01: n11148_o = n10984_o;
      2'b10: n11148_o = n10985_o;
      2'b11: n11148_o = n10986_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11149_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11149_o)
      2'b00: n11150_o = n10987_o;
      2'b01: n11150_o = n10988_o;
      2'b10: n11150_o = n10989_o;
      2'b11: n11150_o = n10990_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11151_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11151_o)
      2'b00: n11152_o = n10991_o;
      2'b01: n11152_o = n10992_o;
      2'b10: n11152_o = n10993_o;
      2'b11: n11152_o = n10994_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11153_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11153_o)
      2'b00: n11154_o = n10995_o;
      2'b01: n11154_o = n10996_o;
      2'b10: n11154_o = n10997_o;
      2'b11: n11154_o = n10998_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11155_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11155_o)
      2'b00: n11156_o = n10999_o;
      2'b01: n11156_o = n11000_o;
      2'b10: n11156_o = n11001_o;
      2'b11: n11156_o = n11002_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11157_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11157_o)
      2'b00: n11158_o = n11003_o;
      2'b01: n11158_o = n11004_o;
      2'b10: n11158_o = n11005_o;
      2'b11: n11158_o = n11006_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11159_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11159_o)
      2'b00: n11160_o = n11007_o;
      2'b01: n11160_o = n11008_o;
      2'b10: n11160_o = n11009_o;
      2'b11: n11160_o = n11010_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11161_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11161_o)
      2'b00: n11162_o = n11011_o;
      2'b01: n11162_o = n11012_o;
      2'b10: n11162_o = n11013_o;
      2'b11: n11162_o = n11014_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11163_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11163_o)
      2'b00: n11164_o = n11015_o;
      2'b01: n11164_o = n11016_o;
      2'b10: n11164_o = n11017_o;
      2'b11: n11164_o = n11018_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11165_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11165_o)
      2'b00: n11166_o = n11019_o;
      2'b01: n11166_o = n11020_o;
      2'b10: n11166_o = n11021_o;
      2'b11: n11166_o = n11022_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11167_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11167_o)
      2'b00: n11168_o = n11023_o;
      2'b01: n11168_o = n11024_o;
      2'b10: n11168_o = n11025_o;
      2'b11: n11168_o = n11026_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11169_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11169_o)
      2'b00: n11170_o = n11027_o;
      2'b01: n11170_o = n11028_o;
      2'b10: n11170_o = n11029_o;
      2'b11: n11170_o = n11030_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11171_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11171_o)
      2'b00: n11172_o = n11031_o;
      2'b01: n11172_o = n11032_o;
      2'b10: n11172_o = n11033_o;
      2'b11: n11172_o = n11034_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11173_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11173_o)
      2'b00: n11174_o = n11035_o;
      2'b01: n11174_o = n11036_o;
      2'b10: n11174_o = n11037_o;
      2'b11: n11174_o = n11038_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11175_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11175_o)
      2'b00: n11176_o = n11039_o;
      2'b01: n11176_o = n11040_o;
      2'b10: n11176_o = n11041_o;
      2'b11: n11176_o = n11042_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11177_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11177_o)
      2'b00: n11178_o = n11043_o;
      2'b01: n11178_o = n11044_o;
      2'b10: n11178_o = n11045_o;
      2'b11: n11178_o = n11046_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11179_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11179_o)
      2'b00: n11180_o = n11047_o;
      2'b01: n11180_o = n11048_o;
      2'b10: n11180_o = n11049_o;
      2'b11: n11180_o = n11050_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11181_o = n9748_o[1:0];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11181_o)
      2'b00: n11182_o = n11051_o;
      2'b01: n11182_o = n11052_o;
      2'b10: n11182_o = n11053_o;
      2'b11: n11182_o = n11054_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11183_o = n9748_o[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11183_o)
      2'b00: n11184_o = n11056_o;
      2'b01: n11184_o = n11058_o;
      2'b10: n11184_o = n11060_o;
      2'b11: n11184_o = n11062_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11185_o = n9748_o[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11185_o)
      2'b00: n11186_o = n11064_o;
      2'b01: n11186_o = n11066_o;
      2'b10: n11186_o = n11068_o;
      2'b11: n11186_o = n11070_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11187_o = n9748_o[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11187_o)
      2'b00: n11188_o = n11072_o;
      2'b01: n11188_o = n11074_o;
      2'b10: n11188_o = n11076_o;
      2'b11: n11188_o = n11078_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11189_o = n9748_o[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11189_o)
      2'b00: n11190_o = n11080_o;
      2'b01: n11190_o = n11082_o;
      2'b10: n11190_o = n11084_o;
      2'b11: n11190_o = n11086_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11191_o = n9748_o[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11191_o)
      2'b00: n11192_o = n11088_o;
      2'b01: n11192_o = n11090_o;
      2'b10: n11192_o = n11092_o;
      2'b11: n11192_o = n11094_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11193_o = n9748_o[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11193_o)
      2'b00: n11194_o = n11096_o;
      2'b01: n11194_o = n11098_o;
      2'b10: n11194_o = n11100_o;
      2'b11: n11194_o = n11102_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11195_o = n9748_o[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11195_o)
      2'b00: n11196_o = n11104_o;
      2'b01: n11196_o = n11106_o;
      2'b10: n11196_o = n11108_o;
      2'b11: n11196_o = n11110_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11197_o = n9748_o[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11197_o)
      2'b00: n11198_o = n11112_o;
      2'b01: n11198_o = n11114_o;
      2'b10: n11198_o = n11116_o;
      2'b11: n11198_o = n11118_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11199_o = n9748_o[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11199_o)
      2'b00: n11200_o = n11120_o;
      2'b01: n11200_o = n11122_o;
      2'b10: n11200_o = n11124_o;
      2'b11: n11200_o = n11126_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11201_o = n9748_o[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11201_o)
      2'b00: n11202_o = n11128_o;
      2'b01: n11202_o = n11130_o;
      2'b10: n11202_o = n11132_o;
      2'b11: n11202_o = n11134_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11203_o = n9748_o[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11203_o)
      2'b00: n11204_o = n11136_o;
      2'b01: n11204_o = n11138_o;
      2'b10: n11204_o = n11140_o;
      2'b11: n11204_o = n11142_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11205_o = n9748_o[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11205_o)
      2'b00: n11206_o = n11144_o;
      2'b01: n11206_o = n11146_o;
      2'b10: n11206_o = n11148_o;
      2'b11: n11206_o = n11150_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11207_o = n9748_o[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11207_o)
      2'b00: n11208_o = n11152_o;
      2'b01: n11208_o = n11154_o;
      2'b10: n11208_o = n11156_o;
      2'b11: n11208_o = n11158_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11209_o = n9748_o[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11209_o)
      2'b00: n11210_o = n11160_o;
      2'b01: n11210_o = n11162_o;
      2'b10: n11210_o = n11164_o;
      2'b11: n11210_o = n11166_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11211_o = n9748_o[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11211_o)
      2'b00: n11212_o = n11168_o;
      2'b01: n11212_o = n11170_o;
      2'b10: n11212_o = n11172_o;
      2'b11: n11212_o = n11174_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11213_o = n9748_o[3:2];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11213_o)
      2'b00: n11214_o = n11176_o;
      2'b01: n11214_o = n11178_o;
      2'b10: n11214_o = n11180_o;
      2'b11: n11214_o = n11182_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11215_o = n9748_o[5:4];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11215_o)
      2'b00: n11216_o = n11184_o;
      2'b01: n11216_o = n11186_o;
      2'b10: n11216_o = n11188_o;
      2'b11: n11216_o = n11190_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11217_o = n9748_o[5:4];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11217_o)
      2'b00: n11218_o = n11192_o;
      2'b01: n11218_o = n11194_o;
      2'b10: n11218_o = n11196_o;
      2'b11: n11218_o = n11198_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11219_o = n9748_o[5:4];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11219_o)
      2'b00: n11220_o = n11200_o;
      2'b01: n11220_o = n11202_o;
      2'b10: n11220_o = n11204_o;
      2'b11: n11220_o = n11206_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11221_o = n9748_o[5:4];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11221_o)
      2'b00: n11222_o = n11208_o;
      2'b01: n11222_o = n11210_o;
      2'b10: n11222_o = n11212_o;
      2'b11: n11222_o = n11214_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  assign n11223_o = n9748_o[7:6];
  /* ../neorv32/rtl/core/neorv32_fifo.vhd:227:31  */
  always @*
    case (n11223_o)
      2'b00: n11224_o = n11216_o;
      2'b01: n11224_o = n11218_o;
      2'b10: n11224_o = n11220_o;
      2'b11: n11224_o = n11222_o;
    endcase
endmodule

module neorv32_cpu_bus_32_0_4
  (input  clk_i,
   input  rstn_i,
   input  ctrl_i_rf_wb_en,
   input  [4:0] ctrl_i_rf_rs1,
   input  [4:0] ctrl_i_rf_rs2,
   input  [4:0] ctrl_i_rf_rs3,
   input  [4:0] ctrl_i_rf_rd,
   input  [1:0] ctrl_i_rf_mux,
   input  ctrl_i_rf_zero_we,
   input  [2:0] ctrl_i_alu_op,
   input  ctrl_i_alu_opa_mux,
   input  ctrl_i_alu_opb_mux,
   input  ctrl_i_alu_unsigned,
   input  [2:0] ctrl_i_alu_frm,
   input  [5:0] ctrl_i_alu_cp_trig,
   input  ctrl_i_bus_req,
   input  ctrl_i_bus_mo_we,
   input  ctrl_i_bus_fence,
   input  ctrl_i_bus_fencei,
   input  ctrl_i_bus_priv,
   input  [2:0] ctrl_i_ir_funct3,
   input  [11:0] ctrl_i_ir_funct12,
   input  [6:0] ctrl_i_ir_opcode,
   input  ctrl_i_cpu_priv,
   input  ctrl_i_cpu_sleep,
   input  ctrl_i_cpu_trap,
   input  ctrl_i_cpu_debug,
   input  [31:0] fetch_pc_i,
   input  [31:0] addr_i,
   input  [31:0] wdata_i,
   input  [543:0] pmp_addr_i,
   input  [127:0] pmp_ctrl_i,
   input  [31:0] d_bus_rdata_i,
   input  d_bus_ack_i,
   input  d_bus_err_i,
   output i_pmp_fault_o,
   output [31:0] rdata_o,
   output [31:0] mar_o,
   output d_wait_o,
   output ma_load_o,
   output ma_store_o,
   output be_load_o,
   output be_store_o,
   output [31:0] d_bus_addr_o,
   output [31:0] d_bus_wdata_o,
   output [3:0] d_bus_ben_o,
   output d_bus_we_o,
   output d_bus_re_o,
   output d_bus_fence_o,
   output d_bus_priv_o);
  wire [69:0] n9046_o;
  wire data_sign;
  wire [31:0] mar;
  wire misaligned;
  wire [3:0] arbiter;
  wire if_pmp_fault;
  wire ld_pmp_fault;
  wire st_pmp_fault;
  wire n9064_o;
  wire [1:0] n9065_o;
  wire n9067_o;
  wire n9068_o;
  wire n9070_o;
  wire n9071_o;
  wire n9072_o;
  wire n9073_o;
  wire n9075_o;
  wire [2:0] n9076_o;
  reg n9079_o;
  wire n9087_o;
  wire [1:0] n9088_o;
  wire [7:0] n9089_o;
  wire [7:0] n9090_o;
  wire [7:0] n9091_o;
  wire [7:0] n9092_o;
  wire [1:0] n9093_o;
  localparam [3:0] n9096_o = 4'b0000;
  wire n9100_o;
  wire [15:0] n9101_o;
  wire [15:0] n9102_o;
  wire n9103_o;
  wire n9104_o;
  wire [3:0] n9107_o;
  wire n9109_o;
  wire [1:0] n9110_o;
  wire [7:0] n9111_o;
  wire [7:0] n9112_o;
  reg [7:0] n9113_o;
  wire [7:0] n9114_o;
  wire [7:0] n9115_o;
  reg [7:0] n9116_o;
  wire [7:0] n9117_o;
  wire [7:0] n9118_o;
  reg [7:0] n9119_o;
  wire [7:0] n9120_o;
  wire [7:0] n9121_o;
  reg [7:0] n9122_o;
  reg [3:0] n9124_o;
  wire [31:0] n9126_o;
  wire [1:0] n9135_o;
  wire [1:0] n9136_o;
  wire [7:0] n9137_o;
  wire n9138_o;
  wire n9139_o;
  wire n9140_o;
  wire n9141_o;
  wire n9142_o;
  wire n9143_o;
  wire n9144_o;
  wire n9145_o;
  wire n9146_o;
  wire n9147_o;
  wire n9148_o;
  wire n9149_o;
  wire n9150_o;
  wire n9151_o;
  wire n9152_o;
  wire n9153_o;
  wire n9154_o;
  wire n9155_o;
  wire n9156_o;
  wire n9157_o;
  wire n9158_o;
  wire n9159_o;
  wire n9160_o;
  wire n9161_o;
  wire n9162_o;
  wire n9163_o;
  wire n9164_o;
  wire n9165_o;
  wire n9166_o;
  wire n9167_o;
  wire n9168_o;
  wire n9169_o;
  wire n9170_o;
  wire n9171_o;
  wire n9172_o;
  wire n9173_o;
  wire n9174_o;
  wire n9175_o;
  wire n9176_o;
  wire n9177_o;
  wire n9178_o;
  wire n9179_o;
  wire n9180_o;
  wire n9181_o;
  wire n9182_o;
  wire n9183_o;
  wire n9184_o;
  wire n9185_o;
  wire [3:0] n9186_o;
  wire [3:0] n9187_o;
  wire [3:0] n9188_o;
  wire [3:0] n9189_o;
  wire [3:0] n9190_o;
  wire [3:0] n9191_o;
  wire [15:0] n9192_o;
  wire [7:0] n9193_o;
  wire [23:0] n9194_o;
  wire n9196_o;
  wire [7:0] n9197_o;
  wire n9198_o;
  wire n9199_o;
  wire n9200_o;
  wire n9201_o;
  wire n9202_o;
  wire n9203_o;
  wire n9204_o;
  wire n9205_o;
  wire n9206_o;
  wire n9207_o;
  wire n9208_o;
  wire n9209_o;
  wire n9210_o;
  wire n9211_o;
  wire n9212_o;
  wire n9213_o;
  wire n9214_o;
  wire n9215_o;
  wire n9216_o;
  wire n9217_o;
  wire n9218_o;
  wire n9219_o;
  wire n9220_o;
  wire n9221_o;
  wire n9222_o;
  wire n9223_o;
  wire n9224_o;
  wire n9225_o;
  wire n9226_o;
  wire n9227_o;
  wire n9228_o;
  wire n9229_o;
  wire n9230_o;
  wire n9231_o;
  wire n9232_o;
  wire n9233_o;
  wire n9234_o;
  wire n9235_o;
  wire n9236_o;
  wire n9237_o;
  wire n9238_o;
  wire n9239_o;
  wire n9240_o;
  wire n9241_o;
  wire n9242_o;
  wire n9243_o;
  wire n9244_o;
  wire n9245_o;
  wire [3:0] n9246_o;
  wire [3:0] n9247_o;
  wire [3:0] n9248_o;
  wire [3:0] n9249_o;
  wire [3:0] n9250_o;
  wire [3:0] n9251_o;
  wire [15:0] n9252_o;
  wire [7:0] n9253_o;
  wire [23:0] n9254_o;
  wire n9256_o;
  wire [7:0] n9257_o;
  wire n9258_o;
  wire n9259_o;
  wire n9260_o;
  wire n9261_o;
  wire n9262_o;
  wire n9263_o;
  wire n9264_o;
  wire n9265_o;
  wire n9266_o;
  wire n9267_o;
  wire n9268_o;
  wire n9269_o;
  wire n9270_o;
  wire n9271_o;
  wire n9272_o;
  wire n9273_o;
  wire n9274_o;
  wire n9275_o;
  wire n9276_o;
  wire n9277_o;
  wire n9278_o;
  wire n9279_o;
  wire n9280_o;
  wire n9281_o;
  wire n9282_o;
  wire n9283_o;
  wire n9284_o;
  wire n9285_o;
  wire n9286_o;
  wire n9287_o;
  wire n9288_o;
  wire n9289_o;
  wire n9290_o;
  wire n9291_o;
  wire n9292_o;
  wire n9293_o;
  wire n9294_o;
  wire n9295_o;
  wire n9296_o;
  wire n9297_o;
  wire n9298_o;
  wire n9299_o;
  wire n9300_o;
  wire n9301_o;
  wire n9302_o;
  wire n9303_o;
  wire n9304_o;
  wire n9305_o;
  wire [3:0] n9306_o;
  wire [3:0] n9307_o;
  wire [3:0] n9308_o;
  wire [3:0] n9309_o;
  wire [3:0] n9310_o;
  wire [3:0] n9311_o;
  wire [15:0] n9312_o;
  wire [7:0] n9313_o;
  wire [23:0] n9314_o;
  wire n9316_o;
  wire [7:0] n9317_o;
  wire n9318_o;
  wire n9319_o;
  wire n9320_o;
  wire n9321_o;
  wire n9322_o;
  wire n9323_o;
  wire n9324_o;
  wire n9325_o;
  wire n9326_o;
  wire n9327_o;
  wire n9328_o;
  wire n9329_o;
  wire n9330_o;
  wire n9331_o;
  wire n9332_o;
  wire n9333_o;
  wire n9334_o;
  wire n9335_o;
  wire n9336_o;
  wire n9337_o;
  wire n9338_o;
  wire n9339_o;
  wire n9340_o;
  wire n9341_o;
  wire n9342_o;
  wire n9343_o;
  wire n9344_o;
  wire n9345_o;
  wire n9346_o;
  wire n9347_o;
  wire n9348_o;
  wire n9349_o;
  wire n9350_o;
  wire n9351_o;
  wire n9352_o;
  wire n9353_o;
  wire n9354_o;
  wire n9355_o;
  wire n9356_o;
  wire n9357_o;
  wire n9358_o;
  wire n9359_o;
  wire n9360_o;
  wire n9361_o;
  wire n9362_o;
  wire n9363_o;
  wire n9364_o;
  wire n9365_o;
  wire [3:0] n9366_o;
  wire [3:0] n9367_o;
  wire [3:0] n9368_o;
  wire [3:0] n9369_o;
  wire [3:0] n9370_o;
  wire [3:0] n9371_o;
  wire [15:0] n9372_o;
  wire [7:0] n9373_o;
  wire [23:0] n9374_o;
  wire [2:0] n9375_o;
  reg [7:0] n9376_o;
  reg [23:0] n9377_o;
  wire n9379_o;
  wire n9380_o;
  wire n9381_o;
  wire [15:0] n9382_o;
  wire n9383_o;
  wire n9384_o;
  wire n9385_o;
  wire n9386_o;
  wire n9387_o;
  wire n9388_o;
  wire n9389_o;
  wire n9390_o;
  wire n9391_o;
  wire n9392_o;
  wire n9393_o;
  wire n9394_o;
  wire n9395_o;
  wire n9396_o;
  wire n9397_o;
  wire n9398_o;
  wire n9399_o;
  wire n9400_o;
  wire n9401_o;
  wire n9402_o;
  wire n9403_o;
  wire n9404_o;
  wire n9405_o;
  wire n9406_o;
  wire n9407_o;
  wire n9408_o;
  wire n9409_o;
  wire n9410_o;
  wire n9411_o;
  wire n9412_o;
  wire n9413_o;
  wire n9414_o;
  wire [3:0] n9415_o;
  wire [3:0] n9416_o;
  wire [3:0] n9417_o;
  wire [3:0] n9418_o;
  wire [15:0] n9419_o;
  wire [15:0] n9420_o;
  wire n9421_o;
  wire n9422_o;
  wire n9423_o;
  wire n9424_o;
  wire n9425_o;
  wire n9426_o;
  wire n9427_o;
  wire n9428_o;
  wire n9429_o;
  wire n9430_o;
  wire n9431_o;
  wire n9432_o;
  wire n9433_o;
  wire n9434_o;
  wire n9435_o;
  wire n9436_o;
  wire n9437_o;
  wire n9438_o;
  wire n9439_o;
  wire n9440_o;
  wire n9441_o;
  wire n9442_o;
  wire n9443_o;
  wire n9444_o;
  wire n9445_o;
  wire n9446_o;
  wire n9447_o;
  wire n9448_o;
  wire n9449_o;
  wire n9450_o;
  wire n9451_o;
  wire n9452_o;
  wire [3:0] n9453_o;
  wire [3:0] n9454_o;
  wire [3:0] n9455_o;
  wire [3:0] n9456_o;
  wire [15:0] n9457_o;
  wire [31:0] n9458_o;
  wire [31:0] n9459_o;
  wire [31:0] n9460_o;
  wire n9462_o;
  wire [1:0] n9463_o;
  wire [7:0] n9464_o;
  wire [7:0] n9465_o;
  reg [7:0] n9466_o;
  wire [23:0] n9467_o;
  wire [23:0] n9468_o;
  reg [23:0] n9469_o;
  wire [31:0] n9471_o;
  wire n9476_o;
  wire n9477_o;
  wire n9479_o;
  wire n9485_o;
  wire n9486_o;
  wire n9487_o;
  wire n9489_o;
  wire n9490_o;
  wire n9492_o;
  wire n9493_o;
  wire n9494_o;
  wire n9495_o;
  wire n9496_o;
  wire n9497_o;
  wire n9498_o;
  wire n9499_o;
  wire n9500_o;
  wire n9502_o;
  wire n9503_o;
  wire n9504_o;
  wire n9505_o;
  wire n9507_o;
  wire n9508_o;
  wire [1:0] n9509_o;
  wire [1:0] n9510_o;
  wire [1:0] n9511_o;
  wire n9512_o;
  wire [1:0] n9513_o;
  wire [1:0] n9514_o;
  wire [1:0] n9515_o;
  wire [3:0] n9516_o;
  wire [3:0] n9518_o;
  wire n9521_o;
  wire n9523_o;
  wire n9524_o;
  wire n9525_o;
  wire n9526_o;
  wire n9527_o;
  wire n9528_o;
  wire n9531_o;
  wire n9532_o;
  wire n9533_o;
  wire n9534_o;
  wire n9535_o;
  wire n9536_o;
  wire n9537_o;
  wire n9540_o;
  wire n9541_o;
  wire n9542_o;
  wire n9543_o;
  wire n9544_o;
  wire n9547_o;
  wire n9548_o;
  wire n9549_o;
  wire n9550_o;
  wire n9551_o;
  wire n9552_o;
  wire n9554_o;
  wire n9555_o;
  wire n9556_o;
  wire n9557_o;
  wire n9558_o;
  wire n9559_o;
  wire n9560_o;
  wire n9561_o;
  wire n9562_o;
  wire n9563_o;
  wire n9564_o;
  wire n9565_o;
  wire n9566_o;
  wire n9567_o;
  wire n9568_o;
  wire n9569_o;
  wire n9570_o;
  wire n9571_o;
  wire n9572_o;
  wire n9597_o;
  wire n9602_o;
  wire n9607_o;
  wire [31:0] n9609_o;
  reg [31:0] n9610_q;
  wire n9611_o;
  reg n9612_q;
  reg [3:0] n9613_q;
  reg [31:0] n9616_q;
  wire [31:0] n9617_o;
  reg [31:0] n9618_q;
  wire [3:0] n9619_o;
  reg [3:0] n9620_q;
  wire n9622_o;
  wire n9623_o;
  wire n9624_o;
  wire n9625_o;
  wire n9626_o;
  wire n9627_o;
  wire n9628_o;
  wire n9629_o;
  wire n9630_o;
  wire n9631_o;
  wire n9632_o;
  wire n9633_o;
  wire n9634_o;
  wire n9635_o;
  wire n9636_o;
  wire n9637_o;
  wire [3:0] n9638_o;
  assign i_pmp_fault_o = if_pmp_fault;
  assign rdata_o = n9616_q;
  assign mar_o = mar;
  assign d_wait_o = n9521_o;
  assign ma_load_o = n9528_o;
  assign ma_store_o = n9544_o;
  assign be_load_o = n9537_o;
  assign be_store_o = n9552_o;
  assign d_bus_addr_o = mar;
  assign d_bus_wdata_o = n9618_q;
  assign d_bus_ben_o = n9620_q;
  assign d_bus_we_o = n9561_o;
  assign d_bus_re_o = n9570_o;
  assign d_bus_fence_o = n9571_o;
  assign d_bus_priv_o = n9572_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:257:18  */
  assign n9046_o = {ctrl_i_cpu_debug, ctrl_i_cpu_trap, ctrl_i_cpu_sleep, ctrl_i_cpu_priv, ctrl_i_ir_opcode, ctrl_i_ir_funct12, ctrl_i_ir_funct3, ctrl_i_bus_priv, ctrl_i_bus_fencei, ctrl_i_bus_fence, ctrl_i_bus_mo_we, ctrl_i_bus_req, ctrl_i_alu_cp_trig, ctrl_i_alu_frm, ctrl_i_alu_unsigned, ctrl_i_alu_opb_mux, ctrl_i_alu_opa_mux, ctrl_i_alu_op, ctrl_i_rf_zero_we, ctrl_i_rf_mux, ctrl_i_rf_rd, ctrl_i_rf_rs3, ctrl_i_rf_rs2, ctrl_i_rf_rs1, ctrl_i_rf_wb_en};
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:100:10  */
  assign data_sign = n9477_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:101:10  */
  assign mar = n9610_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:102:10  */
  assign misaligned = n9612_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:111:10  */
  assign arbiter = n9613_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:138:10  */
  assign if_pmp_fault = n9597_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:139:10  */
  assign ld_pmp_fault = n9602_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:140:10  */
  assign st_pmp_fault = n9607_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:149:18  */
  assign n9064_o = n9046_o[40];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:151:30  */
  assign n9065_o = n9046_o[45:44];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:152:11  */
  assign n9067_o = n9065_o == 2'b00;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:153:46  */
  assign n9068_o = addr_i[0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:153:11  */
  assign n9070_o = n9065_o == 2'b01;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:154:46  */
  assign n9071_o = addr_i[1];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:154:59  */
  assign n9072_o = addr_i[0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:154:50  */
  assign n9073_o = n9071_o | n9072_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:154:11  */
  assign n9075_o = n9065_o == 2'b10;
  assign n9076_o = {n9075_o, n9070_o, n9067_o};
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:151:9  */
  always @*
    case (n9076_o)
      3'b100: n9079_o = n9073_o;
      3'b010: n9079_o = n9068_o;
      3'b001: n9079_o = 1'b0;
      default: n9079_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:178:20  */
  assign n9087_o = n9046_o[40];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:180:32  */
  assign n9088_o = n9046_o[45:44];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:184:59  */
  assign n9089_o = wdata_i[7:0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:184:59  */
  assign n9090_o = wdata_i[7:0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:184:59  */
  assign n9091_o = wdata_i[7:0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:184:59  */
  assign n9092_o = wdata_i[7:0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:186:53  */
  assign n9093_o = addr_i[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:182:13  */
  assign n9100_o = n9088_o == 2'b00;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:190:62  */
  assign n9101_o = wdata_i[15:0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:190:62  */
  assign n9102_o = wdata_i[15:0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:192:25  */
  assign n9103_o = addr_i[1];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:192:29  */
  assign n9104_o = ~n9103_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:192:15  */
  assign n9107_o = n9104_o ? 4'b0011 : 4'b1100;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:188:13  */
  assign n9109_o = n9088_o == 2'b01;
  assign n9110_o = {n9109_o, n9100_o};
  assign n9111_o = n9101_o[7:0];
  assign n9112_o = wdata_i[7:0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:180:11  */
  always @*
    case (n9110_o)
      2'b10: n9113_o = n9111_o;
      2'b01: n9113_o = n9089_o;
      default: n9113_o = n9112_o;
    endcase
  assign n9114_o = n9101_o[15:8];
  assign n9115_o = wdata_i[15:8];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:180:11  */
  always @*
    case (n9110_o)
      2'b10: n9116_o = n9114_o;
      2'b01: n9116_o = n9090_o;
      default: n9116_o = n9115_o;
    endcase
  assign n9117_o = n9102_o[7:0];
  assign n9118_o = wdata_i[23:16];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:180:11  */
  always @*
    case (n9110_o)
      2'b10: n9119_o = n9117_o;
      2'b01: n9119_o = n9091_o;
      default: n9119_o = n9118_o;
    endcase
  assign n9120_o = n9102_o[15:8];
  assign n9121_o = wdata_i[31:24];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:180:11  */
  always @*
    case (n9110_o)
      2'b10: n9122_o = n9120_o;
      2'b01: n9122_o = n9092_o;
      default: n9122_o = n9121_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:180:11  */
  always @*
    case (n9110_o)
      2'b10: n9124_o = n9107_o;
      2'b01: n9124_o = n9638_o;
      default: n9124_o = 4'b1111;
    endcase
  assign n9126_o = {n9122_o, n9119_o, n9116_o, n9113_o};
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:269:30  */
  assign n9135_o = n9046_o[45:44];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:272:25  */
  assign n9136_o = mar[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:275:53  */
  assign n9137_o = d_bus_rdata_i[7:0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9138_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9139_o = data_sign & n9138_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9140_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9141_o = data_sign & n9140_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9142_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9143_o = data_sign & n9142_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9144_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9145_o = data_sign & n9144_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9146_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9147_o = data_sign & n9146_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9148_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9149_o = data_sign & n9148_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9150_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9151_o = data_sign & n9150_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9152_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9153_o = data_sign & n9152_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9154_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9155_o = data_sign & n9154_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9156_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9157_o = data_sign & n9156_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9158_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9159_o = data_sign & n9158_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9160_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9161_o = data_sign & n9160_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9162_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9163_o = data_sign & n9162_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9164_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9165_o = data_sign & n9164_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9166_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9167_o = data_sign & n9166_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9168_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9169_o = data_sign & n9168_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9170_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9171_o = data_sign & n9170_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9172_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9173_o = data_sign & n9172_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9174_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9175_o = data_sign & n9174_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9176_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9177_o = data_sign & n9176_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9178_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9179_o = data_sign & n9178_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9180_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9181_o = data_sign & n9180_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9182_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9183_o = data_sign & n9182_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:84  */
  assign n9184_o = d_bus_rdata_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:276:67  */
  assign n9185_o = data_sign & n9184_o;
  assign n9186_o = {n9139_o, n9141_o, n9143_o, n9145_o};
  assign n9187_o = {n9147_o, n9149_o, n9151_o, n9153_o};
  assign n9188_o = {n9155_o, n9157_o, n9159_o, n9161_o};
  assign n9189_o = {n9163_o, n9165_o, n9167_o, n9169_o};
  assign n9190_o = {n9171_o, n9173_o, n9175_o, n9177_o};
  assign n9191_o = {n9179_o, n9181_o, n9183_o, n9185_o};
  assign n9192_o = {n9186_o, n9187_o, n9188_o, n9189_o};
  assign n9193_o = {n9190_o, n9191_o};
  assign n9194_o = {n9192_o, n9193_o};
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:274:15  */
  assign n9196_o = n9136_o == 2'b00;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:278:53  */
  assign n9197_o = d_bus_rdata_i[15:8];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9198_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9199_o = data_sign & n9198_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9200_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9201_o = data_sign & n9200_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9202_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9203_o = data_sign & n9202_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9204_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9205_o = data_sign & n9204_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9206_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9207_o = data_sign & n9206_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9208_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9209_o = data_sign & n9208_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9210_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9211_o = data_sign & n9210_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9212_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9213_o = data_sign & n9212_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9214_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9215_o = data_sign & n9214_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9216_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9217_o = data_sign & n9216_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9218_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9219_o = data_sign & n9218_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9220_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9221_o = data_sign & n9220_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9222_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9223_o = data_sign & n9222_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9224_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9225_o = data_sign & n9224_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9226_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9227_o = data_sign & n9226_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9228_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9229_o = data_sign & n9228_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9230_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9231_o = data_sign & n9230_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9232_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9233_o = data_sign & n9232_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9234_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9235_o = data_sign & n9234_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9236_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9237_o = data_sign & n9236_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9238_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9239_o = data_sign & n9238_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9240_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9241_o = data_sign & n9240_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9242_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9243_o = data_sign & n9242_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:84  */
  assign n9244_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:279:67  */
  assign n9245_o = data_sign & n9244_o;
  assign n9246_o = {n9199_o, n9201_o, n9203_o, n9205_o};
  assign n9247_o = {n9207_o, n9209_o, n9211_o, n9213_o};
  assign n9248_o = {n9215_o, n9217_o, n9219_o, n9221_o};
  assign n9249_o = {n9223_o, n9225_o, n9227_o, n9229_o};
  assign n9250_o = {n9231_o, n9233_o, n9235_o, n9237_o};
  assign n9251_o = {n9239_o, n9241_o, n9243_o, n9245_o};
  assign n9252_o = {n9246_o, n9247_o, n9248_o, n9249_o};
  assign n9253_o = {n9250_o, n9251_o};
  assign n9254_o = {n9252_o, n9253_o};
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:277:15  */
  assign n9256_o = n9136_o == 2'b01;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:281:53  */
  assign n9257_o = d_bus_rdata_i[23:16];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9258_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9259_o = data_sign & n9258_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9260_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9261_o = data_sign & n9260_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9262_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9263_o = data_sign & n9262_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9264_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9265_o = data_sign & n9264_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9266_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9267_o = data_sign & n9266_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9268_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9269_o = data_sign & n9268_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9270_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9271_o = data_sign & n9270_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9272_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9273_o = data_sign & n9272_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9274_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9275_o = data_sign & n9274_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9276_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9277_o = data_sign & n9276_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9278_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9279_o = data_sign & n9278_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9280_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9281_o = data_sign & n9280_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9282_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9283_o = data_sign & n9282_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9284_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9285_o = data_sign & n9284_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9286_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9287_o = data_sign & n9286_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9288_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9289_o = data_sign & n9288_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9290_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9291_o = data_sign & n9290_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9292_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9293_o = data_sign & n9292_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9294_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9295_o = data_sign & n9294_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9296_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9297_o = data_sign & n9296_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9298_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9299_o = data_sign & n9298_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9300_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9301_o = data_sign & n9300_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9302_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9303_o = data_sign & n9302_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:84  */
  assign n9304_o = d_bus_rdata_i[23];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:282:67  */
  assign n9305_o = data_sign & n9304_o;
  assign n9306_o = {n9259_o, n9261_o, n9263_o, n9265_o};
  assign n9307_o = {n9267_o, n9269_o, n9271_o, n9273_o};
  assign n9308_o = {n9275_o, n9277_o, n9279_o, n9281_o};
  assign n9309_o = {n9283_o, n9285_o, n9287_o, n9289_o};
  assign n9310_o = {n9291_o, n9293_o, n9295_o, n9297_o};
  assign n9311_o = {n9299_o, n9301_o, n9303_o, n9305_o};
  assign n9312_o = {n9306_o, n9307_o, n9308_o, n9309_o};
  assign n9313_o = {n9310_o, n9311_o};
  assign n9314_o = {n9312_o, n9313_o};
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:280:15  */
  assign n9316_o = n9136_o == 2'b10;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:284:53  */
  assign n9317_o = d_bus_rdata_i[31:24];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9318_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9319_o = data_sign & n9318_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9320_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9321_o = data_sign & n9320_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9322_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9323_o = data_sign & n9322_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9324_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9325_o = data_sign & n9324_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9326_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9327_o = data_sign & n9326_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9328_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9329_o = data_sign & n9328_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9330_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9331_o = data_sign & n9330_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9332_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9333_o = data_sign & n9332_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9334_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9335_o = data_sign & n9334_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9336_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9337_o = data_sign & n9336_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9338_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9339_o = data_sign & n9338_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9340_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9341_o = data_sign & n9340_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9342_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9343_o = data_sign & n9342_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9344_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9345_o = data_sign & n9344_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9346_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9347_o = data_sign & n9346_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9348_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9349_o = data_sign & n9348_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9350_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9351_o = data_sign & n9350_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9352_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9353_o = data_sign & n9352_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9354_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9355_o = data_sign & n9354_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9356_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9357_o = data_sign & n9356_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9358_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9359_o = data_sign & n9358_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9360_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9361_o = data_sign & n9360_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9362_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9363_o = data_sign & n9362_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:84  */
  assign n9364_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:285:67  */
  assign n9365_o = data_sign & n9364_o;
  assign n9366_o = {n9319_o, n9321_o, n9323_o, n9325_o};
  assign n9367_o = {n9327_o, n9329_o, n9331_o, n9333_o};
  assign n9368_o = {n9335_o, n9337_o, n9339_o, n9341_o};
  assign n9369_o = {n9343_o, n9345_o, n9347_o, n9349_o};
  assign n9370_o = {n9351_o, n9353_o, n9355_o, n9357_o};
  assign n9371_o = {n9359_o, n9361_o, n9363_o, n9365_o};
  assign n9372_o = {n9366_o, n9367_o, n9368_o, n9369_o};
  assign n9373_o = {n9370_o, n9371_o};
  assign n9374_o = {n9372_o, n9373_o};
  assign n9375_o = {n9316_o, n9256_o, n9196_o};
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:273:13  */
  always @*
    case (n9375_o)
      3'b100: n9376_o = n9257_o;
      3'b010: n9376_o = n9197_o;
      3'b001: n9376_o = n9137_o;
      default: n9376_o = n9317_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:273:13  */
  always @*
    case (n9375_o)
      3'b100: n9377_o = n9314_o;
      3'b010: n9377_o = n9254_o;
      3'b001: n9377_o = n9194_o;
      default: n9377_o = n9374_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:271:11  */
  assign n9379_o = n9135_o == 2'b00;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:289:20  */
  assign n9380_o = mar[1];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:289:24  */
  assign n9381_o = ~n9380_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:290:52  */
  assign n9382_o = d_bus_rdata_i[15:0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:83  */
  assign n9383_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:66  */
  assign n9384_o = data_sign & n9383_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:83  */
  assign n9385_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:66  */
  assign n9386_o = data_sign & n9385_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:83  */
  assign n9387_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:66  */
  assign n9388_o = data_sign & n9387_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:83  */
  assign n9389_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:66  */
  assign n9390_o = data_sign & n9389_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:83  */
  assign n9391_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:66  */
  assign n9392_o = data_sign & n9391_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:83  */
  assign n9393_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:66  */
  assign n9394_o = data_sign & n9393_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:83  */
  assign n9395_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:66  */
  assign n9396_o = data_sign & n9395_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:83  */
  assign n9397_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:66  */
  assign n9398_o = data_sign & n9397_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:83  */
  assign n9399_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:66  */
  assign n9400_o = data_sign & n9399_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:83  */
  assign n9401_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:66  */
  assign n9402_o = data_sign & n9401_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:83  */
  assign n9403_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:66  */
  assign n9404_o = data_sign & n9403_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:83  */
  assign n9405_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:66  */
  assign n9406_o = data_sign & n9405_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:83  */
  assign n9407_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:66  */
  assign n9408_o = data_sign & n9407_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:83  */
  assign n9409_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:66  */
  assign n9410_o = data_sign & n9409_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:83  */
  assign n9411_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:66  */
  assign n9412_o = data_sign & n9411_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:83  */
  assign n9413_o = d_bus_rdata_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:291:66  */
  assign n9414_o = data_sign & n9413_o;
  assign n9415_o = {n9384_o, n9386_o, n9388_o, n9390_o};
  assign n9416_o = {n9392_o, n9394_o, n9396_o, n9398_o};
  assign n9417_o = {n9400_o, n9402_o, n9404_o, n9406_o};
  assign n9418_o = {n9408_o, n9410_o, n9412_o, n9414_o};
  assign n9419_o = {n9415_o, n9416_o, n9417_o, n9418_o};
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:293:52  */
  assign n9420_o = d_bus_rdata_i[31:16];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:83  */
  assign n9421_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:66  */
  assign n9422_o = data_sign & n9421_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:83  */
  assign n9423_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:66  */
  assign n9424_o = data_sign & n9423_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:83  */
  assign n9425_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:66  */
  assign n9426_o = data_sign & n9425_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:83  */
  assign n9427_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:66  */
  assign n9428_o = data_sign & n9427_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:83  */
  assign n9429_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:66  */
  assign n9430_o = data_sign & n9429_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:83  */
  assign n9431_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:66  */
  assign n9432_o = data_sign & n9431_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:83  */
  assign n9433_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:66  */
  assign n9434_o = data_sign & n9433_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:83  */
  assign n9435_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:66  */
  assign n9436_o = data_sign & n9435_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:83  */
  assign n9437_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:66  */
  assign n9438_o = data_sign & n9437_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:83  */
  assign n9439_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:66  */
  assign n9440_o = data_sign & n9439_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:83  */
  assign n9441_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:66  */
  assign n9442_o = data_sign & n9441_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:83  */
  assign n9443_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:66  */
  assign n9444_o = data_sign & n9443_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:83  */
  assign n9445_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:66  */
  assign n9446_o = data_sign & n9445_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:83  */
  assign n9447_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:66  */
  assign n9448_o = data_sign & n9447_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:83  */
  assign n9449_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:66  */
  assign n9450_o = data_sign & n9449_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:83  */
  assign n9451_o = d_bus_rdata_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:294:66  */
  assign n9452_o = data_sign & n9451_o;
  assign n9453_o = {n9422_o, n9424_o, n9426_o, n9428_o};
  assign n9454_o = {n9430_o, n9432_o, n9434_o, n9436_o};
  assign n9455_o = {n9438_o, n9440_o, n9442_o, n9444_o};
  assign n9456_o = {n9446_o, n9448_o, n9450_o, n9452_o};
  assign n9457_o = {n9453_o, n9454_o, n9455_o, n9456_o};
  assign n9458_o = {n9457_o, n9420_o};
  assign n9459_o = {n9419_o, n9382_o};
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:289:13  */
  assign n9460_o = n9381_o ? n9459_o : n9458_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:288:11  */
  assign n9462_o = n9135_o == 2'b01;
  assign n9463_o = {n9462_o, n9379_o};
  assign n9464_o = n9460_o[7:0];
  assign n9465_o = d_bus_rdata_i[7:0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:269:9  */
  always @*
    case (n9463_o)
      2'b10: n9466_o = n9464_o;
      2'b01: n9466_o = n9376_o;
      default: n9466_o = n9465_o;
    endcase
  assign n9467_o = n9460_o[31:8];
  assign n9468_o = d_bus_rdata_i[31:8];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:269:9  */
  always @*
    case (n9463_o)
      2'b10: n9469_o = n9467_o;
      2'b01: n9469_o = n9377_o;
      default: n9469_o = n9468_o;
    endcase
  assign n9471_o = {n9469_o, n9466_o};
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:378:36  */
  assign n9476_o = n9046_o[46];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:378:16  */
  assign n9477_o = ~n9476_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:385:16  */
  assign n9479_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:392:19  */
  assign n9485_o = arbiter[0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:392:24  */
  assign n9486_o = ~n9485_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:393:20  */
  assign n9487_o = n9046_o[39];
  assign n9489_o = arbiter[0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:393:9  */
  assign n9490_o = n9487_o ? 1'b1 : n9489_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:400:30  */
  assign n9492_o = n9046_o[64];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:400:54  */
  assign n9493_o = arbiter[3];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:400:41  */
  assign n9494_o = n9492_o & n9493_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:399:32  */
  assign n9495_o = d_bus_err_i | n9494_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:401:30  */
  assign n9496_o = n9046_o[64];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:401:34  */
  assign n9497_o = ~n9496_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:401:54  */
  assign n9498_o = arbiter[2];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:401:41  */
  assign n9499_o = n9497_o & n9498_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:400:72  */
  assign n9500_o = n9495_o | n9499_o;
  assign n9502_o = arbiter[1];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:399:9  */
  assign n9503_o = n9500_o ? 1'b1 : n9502_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:405:43  */
  assign n9504_o = n9046_o[68];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:405:32  */
  assign n9505_o = d_bus_ack_i | n9504_o;
  assign n9507_o = arbiter[0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:405:9  */
  assign n9508_o = n9505_o ? 1'b0 : n9507_o;
  assign n9509_o = {n9503_o, n9508_o};
  assign n9510_o = {1'b0, n9490_o};
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:392:7  */
  assign n9511_o = n9486_o ? n9510_o : n9509_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:410:18  */
  assign n9512_o = n9046_o[40];
  assign n9513_o = {st_pmp_fault, ld_pmp_fault};
  assign n9514_o = arbiter[3:2];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:410:7  */
  assign n9515_o = n9512_o ? n9513_o : n9514_o;
  assign n9516_o = {n9515_o, n9511_o};
  assign n9518_o = {1'b0, 1'b0, 1'b0, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:418:15  */
  assign n9521_o = ~d_bus_ack_i;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:421:35  */
  assign n9523_o = arbiter[0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:421:68  */
  assign n9524_o = n9046_o[64];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:421:72  */
  assign n9525_o = ~n9524_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:421:47  */
  assign n9526_o = n9523_o & n9525_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:421:79  */
  assign n9527_o = n9526_o & misaligned;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:421:21  */
  assign n9528_o = n9527_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:422:35  */
  assign n9531_o = arbiter[0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:422:68  */
  assign n9532_o = n9046_o[64];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:422:72  */
  assign n9533_o = ~n9532_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:422:47  */
  assign n9534_o = n9531_o & n9533_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:422:92  */
  assign n9535_o = arbiter[1];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:422:79  */
  assign n9536_o = n9534_o & n9535_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:422:21  */
  assign n9537_o = n9536_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:423:35  */
  assign n9540_o = arbiter[0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:423:68  */
  assign n9541_o = n9046_o[64];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:423:47  */
  assign n9542_o = n9540_o & n9541_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:423:79  */
  assign n9543_o = n9542_o & misaligned;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:423:21  */
  assign n9544_o = n9543_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:424:35  */
  assign n9547_o = arbiter[0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:424:68  */
  assign n9548_o = n9046_o[64];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:424:47  */
  assign n9549_o = n9547_o & n9548_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:424:92  */
  assign n9550_o = arbiter[1];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:424:79  */
  assign n9551_o = n9549_o & n9550_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:424:21  */
  assign n9552_o = n9551_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:427:27  */
  assign n9554_o = n9046_o[39];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:427:60  */
  assign n9555_o = n9046_o[64];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:427:35  */
  assign n9556_o = n9554_o & n9555_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:427:70  */
  assign n9557_o = ~misaligned;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:427:65  */
  assign n9558_o = n9556_o & n9557_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:427:103  */
  assign n9559_o = arbiter[3];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:427:91  */
  assign n9560_o = ~n9559_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:427:86  */
  assign n9561_o = n9558_o & n9560_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:428:27  */
  assign n9562_o = n9046_o[39];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:428:60  */
  assign n9563_o = n9046_o[64];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:428:40  */
  assign n9564_o = ~n9563_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:428:35  */
  assign n9565_o = n9562_o & n9564_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:428:70  */
  assign n9566_o = ~misaligned;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:428:65  */
  assign n9567_o = n9565_o & n9566_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:428:103  */
  assign n9568_o = arbiter[2];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:428:91  */
  assign n9569_o = ~n9568_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:428:86  */
  assign n9570_o = n9567_o & n9569_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:429:27  */
  assign n9571_o = n9046_o[41];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:430:27  */
  assign n9572_o = n9046_o[43];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:535:23  */
  assign n9597_o = 1'b0 ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:536:23  */
  assign n9602_o = 1'b0 ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:537:23  */
  assign n9607_o = 1'b0 ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:148:5  */
  assign n9609_o = n9064_o ? addr_i : mar;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:148:5  */
  always @(posedge clk_i)
    n9610_q <= n9609_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:148:5  */
  assign n9611_o = n9064_o ? n9079_o : misaligned;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:148:5  */
  always @(posedge clk_i)
    n9612_q <= n9611_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:390:5  */
  always @(posedge clk_i or posedge n9479_o)
    if (n9479_o)
      n9613_q <= n9518_o;
    else
      n9613_q <= n9516_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:268:7  */
  always @(posedge clk_i)
    n9616_q <= n9471_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:177:7  */
  assign n9617_o = n9087_o ? n9126_o : n9618_q;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:177:7  */
  always @(posedge clk_i)
    n9618_q <= n9617_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:177:7  */
  assign n9619_o = n9087_o ? n9124_o : n9620_q;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:177:7  */
  always @(posedge clk_i)
    n9620_q <= n9619_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:186:15  */
  assign n9622_o = n9093_o[1];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:186:15  */
  assign n9623_o = ~n9622_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:186:15  */
  assign n9624_o = n9093_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:186:15  */
  assign n9625_o = ~n9624_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:186:15  */
  assign n9626_o = n9623_o & n9625_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:186:15  */
  assign n9627_o = n9623_o & n9624_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:186:15  */
  assign n9628_o = n9622_o & n9625_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:186:15  */
  assign n9629_o = n9622_o & n9624_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:66:5  */
  assign n9630_o = n9096_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:186:15  */
  assign n9631_o = n9626_o ? 1'b1 : n9630_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:64:5  */
  assign n9632_o = n9096_o[1];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:186:15  */
  assign n9633_o = n9627_o ? 1'b1 : n9632_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:62:5  */
  assign n9634_o = n9096_o[2];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:186:15  */
  assign n9635_o = n9628_o ? 1'b1 : n9634_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:57:5  */
  assign n9636_o = n9096_o[3];
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:186:15  */
  assign n9637_o = n9629_o ? 1'b1 : n9636_o;
  /* ../neorv32/rtl/core/neorv32_cpu_bus.vhd:148:5  */
  assign n9638_o = {n9637_o, n9635_o, n9633_o, n9631_o};
endmodule

module neorv32_cpu_alu_32_5e99b7dbd159708117122aa5c1c1bfccec006ed0
  (input  clk_i,
   input  rstn_i,
   input  ctrl_i_rf_wb_en,
   input  [4:0] ctrl_i_rf_rs1,
   input  [4:0] ctrl_i_rf_rs2,
   input  [4:0] ctrl_i_rf_rs3,
   input  [4:0] ctrl_i_rf_rd,
   input  [1:0] ctrl_i_rf_mux,
   input  ctrl_i_rf_zero_we,
   input  [2:0] ctrl_i_alu_op,
   input  ctrl_i_alu_opa_mux,
   input  ctrl_i_alu_opb_mux,
   input  ctrl_i_alu_unsigned,
   input  [2:0] ctrl_i_alu_frm,
   input  [5:0] ctrl_i_alu_cp_trig,
   input  ctrl_i_bus_req,
   input  ctrl_i_bus_mo_we,
   input  ctrl_i_bus_fence,
   input  ctrl_i_bus_fencei,
   input  ctrl_i_bus_priv,
   input  [2:0] ctrl_i_ir_funct3,
   input  [11:0] ctrl_i_ir_funct12,
   input  [6:0] ctrl_i_ir_opcode,
   input  ctrl_i_cpu_priv,
   input  ctrl_i_cpu_sleep,
   input  ctrl_i_cpu_trap,
   input  ctrl_i_cpu_debug,
   input  [31:0] rs1_i,
   input  [31:0] rs2_i,
   input  [31:0] rs3_i,
   input  [31:0] rs4_i,
   input  [31:0] pc_i,
   input  [31:0] imm_i,
   output [1:0] cmp_o,
   output [31:0] res_o,
   output [31:0] add_o,
   output [4:0] fpu_flags_o,
   output exc_o,
   output cp_done_o);
  wire [69:0] n8771_o;
  wire [32:0] cmp_rs1;
  wire [32:0] cmp_rs2;
  wire [1:0] cmp;
  wire [31:0] opa;
  wire [31:0] opb;
  wire [32:0] addsub_res;
  wire [31:0] cp_res;
  wire [10:0] cp_monitor;
  wire [191:0] cp_result;
  wire [5:0] cp_start;
  wire [5:0] cp_valid;
  wire n8778_o;
  wire n8779_o;
  wire n8780_o;
  wire n8781_o;
  wire [32:0] n8782_o;
  wire n8783_o;
  wire n8784_o;
  wire n8785_o;
  wire n8786_o;
  wire [32:0] n8787_o;
  wire n8789_o;
  wire n8790_o;
  wire n8793_o;
  wire n8794_o;
  wire n8796_o;
  wire [31:0] n8797_o;
  wire n8798_o;
  wire [31:0] n8799_o;
  wire n8803_o;
  wire n8804_o;
  wire n8805_o;
  wire n8806_o;
  wire [32:0] n8807_o;
  wire n8808_o;
  wire n8809_o;
  wire n8810_o;
  wire n8811_o;
  wire [32:0] n8812_o;
  wire n8813_o;
  wire [32:0] n8814_o;
  wire [32:0] n8815_o;
  wire [32:0] n8816_o;
  wire [31:0] n8818_o;
  wire [2:0] n8820_o;
  wire [31:0] n8821_o;
  wire n8823_o;
  wire [31:0] n8824_o;
  wire n8826_o;
  wire n8828_o;
  wire n8829_o;
  localparam [31:0] n8830_o = 32'b00000000000000000000000000000000;
  wire [30:0] n8831_o;
  wire n8833_o;
  wire n8835_o;
  wire [31:0] n8836_o;
  wire n8838_o;
  wire [31:0] n8839_o;
  wire n8841_o;
  wire [31:0] n8842_o;
  wire n8844_o;
  wire [31:0] n8845_o;
  wire [7:0] n8846_o;
  wire n8847_o;
  wire n8848_o;
  wire n8849_o;
  wire n8850_o;
  wire n8851_o;
  wire n8852_o;
  wire n8853_o;
  wire n8854_o;
  reg n8855_o;
  wire [30:0] n8856_o;
  wire [30:0] n8857_o;
  wire [30:0] n8858_o;
  wire [30:0] n8859_o;
  wire [30:0] n8860_o;
  wire [30:0] n8861_o;
  wire [30:0] n8862_o;
  wire [30:0] n8863_o;
  reg [30:0] n8864_o;
  wire n8867_o;
  wire n8873_o;
  wire n8874_o;
  wire n8875_o;
  wire n8876_o;
  wire n8877_o;
  wire n8878_o;
  wire n8885_o;
  wire n8887_o;
  wire n8889_o;
  wire n8890_o;
  wire n8891_o;
  wire n8892_o;
  wire n8893_o;
  wire n8894_o;
  wire n8895_o;
  wire n8896_o;
  wire n8897_o;
  wire n8898_o;
  wire n8899_o;
  wire n8900_o;
  wire [5:0] n8903_o;
  wire n8909_o;
  wire n8911_o;
  wire n8913_o;
  wire n8914_o;
  wire n8915_o;
  wire n8916_o;
  wire n8917_o;
  wire n8918_o;
  wire n8919_o;
  wire n8920_o;
  wire n8921_o;
  wire n8922_o;
  wire n8924_o;
  wire n8925_o;
  wire [7:0] n8926_o;
  wire [7:0] n8928_o;
  wire n8929_o;
  wire n8930_o;
  wire n8931_o;
  wire n8933_o;
  wire n8934_o;
  wire n8935_o;
  wire [7:0] n8936_o;
  wire [10:0] n8937_o;
  wire [10:0] n8939_o;
  wire n8942_o;
  wire [5:0] n8943_o;
  wire n8944_o;
  wire n8945_o;
  wire n8946_o;
  wire n8947_o;
  wire n8948_o;
  wire n8949_o;
  wire n8950_o;
  wire n8951_o;
  wire n8952_o;
  wire n8953_o;
  wire n8954_o;
  wire [31:0] n8955_o;
  wire [31:0] n8956_o;
  wire [31:0] n8957_o;
  wire [31:0] n8958_o;
  wire [31:0] n8959_o;
  wire [31:0] n8960_o;
  wire [31:0] n8961_o;
  wire [31:0] n8962_o;
  wire [31:0] n8963_o;
  wire [31:0] n8964_o;
  wire [31:0] n8965_o;
  wire n8966_o;
  wire [4:0] n8968_o;
  wire [31:0] neorv32_cpu_cp_shifter_inst_n8969;
  wire neorv32_cpu_cp_shifter_inst_n8970;
  wire [31:0] neorv32_cpu_cp_shifter_inst_res_o;
  wire neorv32_cpu_cp_shifter_inst_valid_o;
  wire n8971_o;
  wire [4:0] n8972_o;
  wire [4:0] n8973_o;
  wire [4:0] n8974_o;
  wire [4:0] n8975_o;
  wire [1:0] n8976_o;
  wire n8977_o;
  wire [2:0] n8978_o;
  wire n8979_o;
  wire n8980_o;
  wire n8981_o;
  wire [2:0] n8982_o;
  wire [5:0] n8983_o;
  wire n8984_o;
  wire n8985_o;
  wire n8986_o;
  wire n8987_o;
  wire n8988_o;
  wire [2:0] n8989_o;
  wire [11:0] n8990_o;
  wire [6:0] n8991_o;
  wire n8992_o;
  wire n8993_o;
  wire n8994_o;
  wire n8995_o;
  wire n9000_o;
  wire [31:0] neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_n9001;
  wire neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_n9002;
  wire [31:0] neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_res_o;
  wire neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_valid_o;
  wire n9003_o;
  wire [4:0] n9004_o;
  wire [4:0] n9005_o;
  wire [4:0] n9006_o;
  wire [4:0] n9007_o;
  wire [1:0] n9008_o;
  wire n9009_o;
  wire [2:0] n9010_o;
  wire n9011_o;
  wire n9012_o;
  wire n9013_o;
  wire [2:0] n9014_o;
  wire [5:0] n9015_o;
  wire n9016_o;
  wire n9017_o;
  wire n9018_o;
  wire n9019_o;
  wire n9020_o;
  wire [2:0] n9021_o;
  wire [11:0] n9022_o;
  wire [6:0] n9023_o;
  wire n9024_o;
  wire n9025_o;
  wire n9026_o;
  wire n9027_o;
  localparam [4:0] n9035_o = 5'b00000;
  wire [1:0] n9041_o;
  reg [10:0] n9042_q;
  wire [191:0] n9043_o;
  wire [5:0] n9044_o;
  wire [31:0] n9045_o;
  assign cmp_o = cmp;
  assign res_o = n9045_o;
  assign add_o = n8818_o;
  assign fpu_flags_o = n9035_o;
  assign exc_o = n8942_o;
  assign cp_done_o = n8954_o;
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:132:7  */
  assign n8771_o = {ctrl_i_cpu_debug, ctrl_i_cpu_trap, ctrl_i_cpu_sleep, ctrl_i_cpu_priv, ctrl_i_ir_opcode, ctrl_i_ir_funct12, ctrl_i_ir_funct3, ctrl_i_bus_priv, ctrl_i_bus_fencei, ctrl_i_bus_fence, ctrl_i_bus_mo_we, ctrl_i_bus_req, ctrl_i_alu_cp_trig, ctrl_i_alu_frm, ctrl_i_alu_unsigned, ctrl_i_alu_opb_mux, ctrl_i_alu_opa_mux, ctrl_i_alu_op, ctrl_i_rf_zero_we, ctrl_i_rf_mux, ctrl_i_rf_rd, ctrl_i_rf_rs3, ctrl_i_rf_rs2, ctrl_i_rf_rs1, ctrl_i_rf_wb_en};
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:84:10  */
  assign cmp_rs1 = n8782_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:85:10  */
  assign cmp_rs2 = n8787_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:86:10  */
  assign cmp = n9041_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:89:10  */
  assign opa = n8797_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:89:15  */
  assign opb = n8799_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:92:10  */
  assign addsub_res = n8816_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:93:10  */
  assign cp_res = n8965_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:102:10  */
  assign cp_monitor = n9042_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:106:10  */
  assign cp_result = n9043_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:107:10  */
  assign cp_start = n8943_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:108:10  */
  assign cp_valid = n9044_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:114:20  */
  assign n8778_o = rs1_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:114:49  */
  assign n8779_o = n8771_o[29];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:114:38  */
  assign n8780_o = ~n8779_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:114:33  */
  assign n8781_o = n8778_o & n8780_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:114:64  */
  assign n8782_o = {n8781_o, rs1_i};
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:115:20  */
  assign n8783_o = rs2_i[31];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:115:49  */
  assign n8784_o = n8771_o[29];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:115:38  */
  assign n8785_o = ~n8784_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:115:33  */
  assign n8786_o = n8783_o & n8785_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:115:64  */
  assign n8787_o = {n8786_o, rs2_i};
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:117:39  */
  assign n8789_o = rs1_i == rs2_i;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:117:27  */
  assign n8790_o = n8789_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:118:49  */
  assign n8793_o = $signed(cmp_rs1) < $signed(cmp_rs2);
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:118:27  */
  assign n8794_o = n8793_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:124:29  */
  assign n8796_o = n8771_o[27];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:124:16  */
  assign n8797_o = n8796_o ? pc_i : rs1_i;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:125:29  */
  assign n8798_o = n8771_o[28];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:125:16  */
  assign n8799_o = n8798_o ? imm_i : rs2_i;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:134:18  */
  assign n8803_o = opa[31];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:134:45  */
  assign n8804_o = n8771_o[29];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:134:34  */
  assign n8805_o = ~n8804_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:134:29  */
  assign n8806_o = n8803_o & n8805_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:134:60  */
  assign n8807_o = {n8806_o, opa};
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:135:18  */
  assign n8808_o = opb[31];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:135:45  */
  assign n8809_o = n8771_o[29];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:135:34  */
  assign n8810_o = ~n8809_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:135:29  */
  assign n8811_o = n8808_o & n8810_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:135:60  */
  assign n8812_o = {n8811_o, opb};
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:137:22  */
  assign n8813_o = n8771_o[24];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:138:55  */
  assign n8814_o = n8807_o - n8812_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:140:55  */
  assign n8815_o = n8807_o + n8812_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:137:5  */
  assign n8816_o = n8813_o ? n8814_o : n8815_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:145:22  */
  assign n8818_o = addsub_res[31:0];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:152:17  */
  assign n8820_o = n8771_o[26:24];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:153:48  */
  assign n8821_o = addsub_res[31:0];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:153:7  */
  assign n8823_o = n8820_o == 3'b000;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:154:48  */
  assign n8824_o = addsub_res[31:0];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:154:7  */
  assign n8826_o = n8820_o == 3'b001;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:155:7  */
  assign n8828_o = n8820_o == 3'b010;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:156:77  */
  assign n8829_o = addsub_res[32];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:716:26  */
  assign n8831_o = n8830_o[31:1];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:156:7  */
  assign n8833_o = n8820_o == 3'b011;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:157:7  */
  assign n8835_o = n8820_o == 3'b100;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:158:44  */
  assign n8836_o = rs1_i ^ opb;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:158:7  */
  assign n8838_o = n8820_o == 3'b101;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:159:44  */
  assign n8839_o = rs1_i | opb;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:159:7  */
  assign n8841_o = n8820_o == 3'b110;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:160:44  */
  assign n8842_o = rs1_i & opb;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:160:7  */
  assign n8844_o = n8820_o == 3'b111;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:161:48  */
  assign n8845_o = addsub_res[31:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:496:18  */
  assign n8846_o = {n8844_o, n8841_o, n8838_o, n8835_o, n8833_o, n8828_o, n8826_o, n8823_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:484:5  */
  assign n8847_o = n8821_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:496:18  */
  assign n8848_o = n8824_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:464:48  */
  assign n8849_o = cp_res[0];
  assign n8850_o = opb[0];
  assign n8851_o = n8836_o[0];
  assign n8852_o = n8839_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:386:3  */
  assign n8853_o = n8842_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:327:10  */
  assign n8854_o = n8845_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:152:5  */
  always @*
    case (n8846_o)
      8'b10000000: n8855_o = n8853_o;
      8'b01000000: n8855_o = n8852_o;
      8'b00100000: n8855_o = n8851_o;
      8'b00010000: n8855_o = n8850_o;
      8'b00001000: n8855_o = n8829_o;
      8'b00000100: n8855_o = n8849_o;
      8'b00000010: n8855_o = n8848_o;
      8'b00000001: n8855_o = n8847_o;
      default: n8855_o = n8854_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:325:10  */
  assign n8856_o = n8821_o[31:1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:312:10  */
  assign n8857_o = n8824_o[31:1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:311:10  */
  assign n8858_o = cp_res[31:1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:609:5  */
  assign n8859_o = opb[31:1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:7  */
  assign n8860_o = n8836_o[31:1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:7  */
  assign n8861_o = n8839_o[31:1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:7  */
  assign n8862_o = n8842_o[31:1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:7  */
  assign n8863_o = n8845_o[31:1];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:152:5  */
  always @*
    case (n8846_o)
      8'b10000000: n8864_o = n8862_o;
      8'b01000000: n8864_o = n8861_o;
      8'b00100000: n8864_o = n8860_o;
      8'b00010000: n8864_o = n8859_o;
      8'b00001000: n8864_o = n8831_o;
      8'b00000100: n8864_o = n8858_o;
      8'b00000010: n8864_o = n8857_o;
      8'b00000001: n8864_o = n8856_o;
      default: n8864_o = n8863_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:177:16  */
  assign n8867_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:183:36  */
  assign n8873_o = cp_monitor[0];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:183:58  */
  assign n8874_o = cp_monitor[10];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:183:40  */
  assign n8875_o = n8873_o & n8874_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:183:100  */
  assign n8876_o = cp_monitor[1];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:183:85  */
  assign n8877_o = ~n8876_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:183:80  */
  assign n8878_o = n8875_o & n8877_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n8885_o = cp_valid[5];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n8887_o = 1'b0 | n8885_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n8889_o = cp_valid[4];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n8890_o = n8887_o | n8889_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n8891_o = cp_valid[3];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n8892_o = n8890_o | n8891_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n8893_o = cp_valid[2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n8894_o = n8892_o | n8893_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n8895_o = cp_valid[1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n8896_o = n8894_o | n8895_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n8897_o = cp_valid[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n8898_o = n8896_o | n8897_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:185:22  */
  assign n8899_o = cp_monitor[0];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:185:26  */
  assign n8900_o = ~n8899_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:187:32  */
  assign n8903_o = n8771_o[38:33];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n8909_o = n8903_o[5];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n8911_o = 1'b0 | n8909_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n8913_o = n8903_o[4];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n8914_o = n8911_o | n8913_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n8915_o = n8903_o[3];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n8916_o = n8914_o | n8915_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n8917_o = n8903_o[2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n8918_o = n8916_o | n8917_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n8919_o = n8903_o[1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n8920_o = n8918_o | n8919_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n8921_o = n8903_o[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n8922_o = n8920_o | n8921_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:7  */
  assign n8924_o = cp_monitor[0];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:187:9  */
  assign n8925_o = n8922_o ? 1'b1 : n8924_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:191:65  */
  assign n8926_o = cp_monitor[10:3];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:191:70  */
  assign n8928_o = n8926_o + 8'b00000001;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:192:24  */
  assign n8929_o = cp_monitor[1];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:192:46  */
  assign n8930_o = n8771_o[68];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:192:35  */
  assign n8931_o = n8929_o | n8930_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:7  */
  assign n8933_o = cp_monitor[0];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:192:9  */
  assign n8934_o = n8931_o ? 1'b0 : n8933_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:185:7  */
  assign n8935_o = n8900_o ? n8925_o : n8934_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:185:7  */
  assign n8936_o = n8900_o ? 8'b00000000 : n8928_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:7  */
  assign n8937_o = {n8936_o, n8878_o, n8898_o, n8935_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:7  */
  assign n8939_o = {8'b00000000, 1'b0, 1'b0, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:200:23  */
  assign n8942_o = cp_monitor[2];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:204:34  */
  assign n8943_o = n8771_o[38:33];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:208:24  */
  assign n8944_o = cp_valid[0];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:208:39  */
  assign n8945_o = cp_valid[1];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:208:28  */
  assign n8946_o = n8944_o | n8945_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:208:54  */
  assign n8947_o = cp_valid[2];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:208:43  */
  assign n8948_o = n8946_o | n8947_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:208:69  */
  assign n8949_o = cp_valid[3];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:208:58  */
  assign n8950_o = n8948_o | n8949_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:208:84  */
  assign n8951_o = cp_valid[4];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:208:73  */
  assign n8952_o = n8950_o | n8951_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:208:99  */
  assign n8953_o = cp_valid[5];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:208:88  */
  assign n8954_o = n8952_o | n8953_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:212:22  */
  assign n8955_o = cp_result[191:160];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:212:38  */
  assign n8956_o = cp_result[159:128];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:212:26  */
  assign n8957_o = n8955_o | n8956_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:212:54  */
  assign n8958_o = cp_result[127:96];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:212:42  */
  assign n8959_o = n8957_o | n8958_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:212:70  */
  assign n8960_o = cp_result[95:64];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:212:58  */
  assign n8961_o = n8959_o | n8960_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:212:86  */
  assign n8962_o = cp_result[63:32];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:212:74  */
  assign n8963_o = n8961_o | n8962_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:212:102  */
  assign n8964_o = cp_result[31:0];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:212:90  */
  assign n8965_o = n8963_o | n8964_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:227:24  */
  assign n8966_o = cp_start[0];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:230:19  */
  assign n8968_o = opb[4:0];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:232:16  */
  assign neorv32_cpu_cp_shifter_inst_n8969 = neorv32_cpu_cp_shifter_inst_res_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:233:16  */
  assign neorv32_cpu_cp_shifter_inst_n8970 = neorv32_cpu_cp_shifter_inst_valid_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:217:3  */
  neorv32_cpu_cp_shifter_32_5ba93c9db0cff93f52b521d7420e43f6eda2784f neorv32_cpu_cp_shifter_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .ctrl_i_rf_wb_en(n8971_o),
    .ctrl_i_rf_rs1(n8972_o),
    .ctrl_i_rf_rs2(n8973_o),
    .ctrl_i_rf_rs3(n8974_o),
    .ctrl_i_rf_rd(n8975_o),
    .ctrl_i_rf_mux(n8976_o),
    .ctrl_i_rf_zero_we(n8977_o),
    .ctrl_i_alu_op(n8978_o),
    .ctrl_i_alu_opa_mux(n8979_o),
    .ctrl_i_alu_opb_mux(n8980_o),
    .ctrl_i_alu_unsigned(n8981_o),
    .ctrl_i_alu_frm(n8982_o),
    .ctrl_i_alu_cp_trig(n8983_o),
    .ctrl_i_bus_req(n8984_o),
    .ctrl_i_bus_mo_we(n8985_o),
    .ctrl_i_bus_fence(n8986_o),
    .ctrl_i_bus_fencei(n8987_o),
    .ctrl_i_bus_priv(n8988_o),
    .ctrl_i_ir_funct3(n8989_o),
    .ctrl_i_ir_funct12(n8990_o),
    .ctrl_i_ir_opcode(n8991_o),
    .ctrl_i_cpu_priv(n8992_o),
    .ctrl_i_cpu_sleep(n8993_o),
    .ctrl_i_cpu_trap(n8994_o),
    .ctrl_i_cpu_debug(n8995_o),
    .start_i(n8966_o),
    .rs1_i(rs1_i),
    .shamt_i(n8968_o),
    .res_o(neorv32_cpu_cp_shifter_inst_res_o),
    .valid_o(neorv32_cpu_cp_shifter_inst_valid_o));
  assign n8971_o = n8771_o[0];
  assign n8972_o = n8771_o[5:1];
  assign n8973_o = n8771_o[10:6];
  assign n8974_o = n8771_o[15:11];
  assign n8975_o = n8771_o[20:16];
  assign n8976_o = n8771_o[22:21];
  assign n8977_o = n8771_o[23];
  assign n8978_o = n8771_o[26:24];
  assign n8979_o = n8771_o[27];
  assign n8980_o = n8771_o[28];
  assign n8981_o = n8771_o[29];
  assign n8982_o = n8771_o[32:30];
  assign n8983_o = n8771_o[38:33];
  assign n8984_o = n8771_o[39];
  assign n8985_o = n8771_o[40];
  assign n8986_o = n8771_o[41];
  assign n8987_o = n8771_o[42];
  assign n8988_o = n8771_o[43];
  assign n8989_o = n8771_o[46:44];
  assign n8990_o = n8771_o[58:47];
  assign n8991_o = n8771_o[65:59];
  assign n8992_o = n8771_o[66];
  assign n8993_o = n8771_o[67];
  assign n8994_o = n8771_o[68];
  assign n8995_o = n8771_o[69];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:252:26  */
  assign n9000_o = cp_start[1];
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:257:18  */
  assign neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_n9001 = neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_res_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:258:18  */
  assign neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_n9002 = neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_valid_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:241:5  */
  neorv32_cpu_cp_muldiv_32_3f29546453678b855931c174a97d6c0894b8f546 neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .ctrl_i_rf_wb_en(n9003_o),
    .ctrl_i_rf_rs1(n9004_o),
    .ctrl_i_rf_rs2(n9005_o),
    .ctrl_i_rf_rs3(n9006_o),
    .ctrl_i_rf_rd(n9007_o),
    .ctrl_i_rf_mux(n9008_o),
    .ctrl_i_rf_zero_we(n9009_o),
    .ctrl_i_alu_op(n9010_o),
    .ctrl_i_alu_opa_mux(n9011_o),
    .ctrl_i_alu_opb_mux(n9012_o),
    .ctrl_i_alu_unsigned(n9013_o),
    .ctrl_i_alu_frm(n9014_o),
    .ctrl_i_alu_cp_trig(n9015_o),
    .ctrl_i_bus_req(n9016_o),
    .ctrl_i_bus_mo_we(n9017_o),
    .ctrl_i_bus_fence(n9018_o),
    .ctrl_i_bus_fencei(n9019_o),
    .ctrl_i_bus_priv(n9020_o),
    .ctrl_i_ir_funct3(n9021_o),
    .ctrl_i_ir_funct12(n9022_o),
    .ctrl_i_ir_opcode(n9023_o),
    .ctrl_i_cpu_priv(n9024_o),
    .ctrl_i_cpu_sleep(n9025_o),
    .ctrl_i_cpu_trap(n9026_o),
    .ctrl_i_cpu_debug(n9027_o),
    .start_i(n9000_o),
    .rs1_i(rs1_i),
    .rs2_i(rs2_i),
    .res_o(neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_res_o),
    .valid_o(neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_valid_o));
  assign n9003_o = n8771_o[0];
  assign n9004_o = n8771_o[5:1];
  assign n9005_o = n8771_o[10:6];
  assign n9006_o = n8771_o[15:11];
  assign n9007_o = n8771_o[20:16];
  assign n9008_o = n8771_o[22:21];
  assign n9009_o = n8771_o[23];
  assign n9010_o = n8771_o[26:24];
  assign n9011_o = n8771_o[27];
  assign n9012_o = n8771_o[28];
  assign n9013_o = n8771_o[29];
  assign n9014_o = n8771_o[32:30];
  assign n9015_o = n8771_o[38:33];
  assign n9016_o = n8771_o[39];
  assign n9017_o = n8771_o[40];
  assign n9018_o = n8771_o[41];
  assign n9019_o = n8771_o[42];
  assign n9020_o = n8771_o[43];
  assign n9021_o = n8771_o[46:44];
  assign n9022_o = n8771_o[58:47];
  assign n9023_o = n8771_o[65:59];
  assign n9024_o = n8771_o[66];
  assign n9025_o = n8771_o[67];
  assign n9026_o = n8771_o[68];
  assign n9027_o = n8771_o[69];
  assign n9041_o = {n8794_o, n8790_o};
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:182:5  */
  always @(posedge clk_i or posedge n8867_o)
    if (n8867_o)
      n9042_q <= n8939_o;
    else
      n9042_q <= n8937_o;
  /* ../neorv32/rtl/core/neorv32_cpu_alu.vhd:177:5  */
  assign n9043_o = {neorv32_cpu_cp_shifter_inst_n8969, neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_n9001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000};
  assign n9044_o = {1'b0, 1'b0, 1'b0, 1'b0, neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_n9002, neorv32_cpu_cp_shifter_inst_n8970};
  assign n9045_o = {n8864_o, n8855_o};
endmodule

module neorv32_cpu_regfile_32_29e2dcfbb16f63bb0254df7585a15bb6fb5e927d
  (input  clk_i,
   input  ctrl_i_rf_wb_en,
   input  [4:0] ctrl_i_rf_rs1,
   input  [4:0] ctrl_i_rf_rs2,
   input  [4:0] ctrl_i_rf_rs3,
   input  [4:0] ctrl_i_rf_rd,
   input  [1:0] ctrl_i_rf_mux,
   input  ctrl_i_rf_zero_we,
   input  [2:0] ctrl_i_alu_op,
   input  ctrl_i_alu_opa_mux,
   input  ctrl_i_alu_opb_mux,
   input  ctrl_i_alu_unsigned,
   input  [2:0] ctrl_i_alu_frm,
   input  [5:0] ctrl_i_alu_cp_trig,
   input  ctrl_i_bus_req,
   input  ctrl_i_bus_mo_we,
   input  ctrl_i_bus_fence,
   input  ctrl_i_bus_fencei,
   input  ctrl_i_bus_priv,
   input  [2:0] ctrl_i_ir_funct3,
   input  [11:0] ctrl_i_ir_funct12,
   input  [6:0] ctrl_i_ir_opcode,
   input  ctrl_i_cpu_priv,
   input  ctrl_i_cpu_sleep,
   input  ctrl_i_cpu_trap,
   input  ctrl_i_cpu_debug,
   input  [31:0] alu_i,
   input  [31:0] mem_i,
   input  [31:0] csr_i,
   input  [31:0] pc2_i,
   output [31:0] rs1_o,
   output [31:0] rs2_o,
   output [31:0] rs3_o,
   output [31:0] rs4_o);
  wire [69:0] n8698_o;
  wire [31:0] rf_wdata;
  wire rf_we;
  wire rd_zero;
  wire [4:0] opa_addr;
  wire [4:0] opb_addr;
  wire [1:0] n8704_o;
  wire n8706_o;
  wire n8708_o;
  wire n8710_o;
  wire n8712_o;
  wire [3:0] n8713_o;
  reg [31:0] n8714_o;
  wire n8717_o;
  wire [4:0] n8718_o;
  wire [4:0] n8719_o;
  wire n8720_o;
  wire [4:0] n8721_o;
  wire [4:0] n8722_o;
  wire [4:0] n8723_o;
  wire [4:0] n8729_o;
  wire n8731_o;
  wire n8732_o;
  wire n8734_o;
  wire n8735_o;
  wire n8736_o;
  wire n8737_o;
  wire n8738_o;
  reg [31:0] n8764_q;
  reg [31:0] n8765_q;
  reg [31:0] n8767_data; // mem_rd
  reg [31:0] n8769_data; // mem_rd
  assign rs1_o = n8769_data;
  assign rs2_o = n8767_data;
  assign rs3_o = n8764_q;
  assign rs4_o = n8765_q;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8698_o = {ctrl_i_cpu_debug, ctrl_i_cpu_trap, ctrl_i_cpu_sleep, ctrl_i_cpu_priv, ctrl_i_ir_opcode, ctrl_i_ir_funct12, ctrl_i_ir_funct3, ctrl_i_bus_priv, ctrl_i_bus_fencei, ctrl_i_bus_fence, ctrl_i_bus_mo_we, ctrl_i_bus_req, ctrl_i_alu_cp_trig, ctrl_i_alu_frm, ctrl_i_alu_unsigned, ctrl_i_alu_opb_mux, ctrl_i_alu_opa_mux, ctrl_i_alu_op, ctrl_i_rf_zero_we, ctrl_i_rf_mux, ctrl_i_rf_rd, ctrl_i_rf_rs3, ctrl_i_rf_rs2, ctrl_i_rf_rs1, ctrl_i_rf_wb_en};
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:87:10  */
  assign rf_wdata = n8714_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:88:10  */
  assign rf_we = n8738_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:89:10  */
  assign rd_zero = n8732_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:136:55  */
  assign opa_addr = n8718_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:137:55  */
  assign opb_addr = n8723_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:101:17  */
  assign n8704_o = n8698_o[22:21];
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:102:7  */
  assign n8706_o = n8704_o == 2'b00;
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:103:7  */
  assign n8708_o = n8704_o == 2'b01;
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:104:7  */
  assign n8710_o = n8704_o == 2'b10;
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:105:7  */
  assign n8712_o = n8704_o == 2'b11;
  assign n8713_o = {n8712_o, n8710_o, n8708_o, n8706_o};
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:101:5  */
  always @*
    case (n8713_o)
      4'b1000: n8714_o = pc2_i;
      4'b0100: n8714_o = csr_i;
      4'b0010: n8714_o = mem_i;
      4'b0001: n8714_o = alu_i;
      default: n8714_o = alu_i;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:114:36  */
  assign n8717_o = n8698_o[23];
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:114:23  */
  assign n8718_o = n8717_o ? 5'b00000 : n8721_o;
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:115:22  */
  assign n8719_o = n8698_o[20:16];
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:115:41  */
  assign n8720_o = n8698_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:114:54  */
  assign n8721_o = n8720_o ? n8719_o : n8722_o;
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:116:22  */
  assign n8722_o = n8698_o[5:1];
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:117:22  */
  assign n8723_o = n8698_o[10:6];
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:122:31  */
  assign n8729_o = n8698_o[20:16];
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:122:37  */
  assign n8731_o = n8729_o == 5'b00000;
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:122:18  */
  assign n8732_o = n8731_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:123:22  */
  assign n8734_o = n8698_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:123:36  */
  assign n8735_o = ~rd_zero;
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:123:31  */
  assign n8736_o = n8734_o & n8735_o;
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:123:60  */
  assign n8737_o = n8698_o[23];
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:123:50  */
  assign n8738_o = n8736_o | n8737_o;
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:132:7  */
  always @(posedge clk_i)
    n8764_q <= 32'b00000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:132:7  */
  always @(posedge clk_i)
    n8765_q <= 32'b00000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:74:5  */
  reg [31:0] reg_file[31:0] ; // memory
  always @(posedge clk_i)
    if (1'b1)
      n8767_data <= reg_file[opb_addr];
  always @(posedge clk_i)
    if (1'b1)
      n8769_data <= reg_file[opa_addr];
  always @(posedge clk_i)
    if (rf_we)
      reg_file[opa_addr] <= rf_wdata;
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:73:5  */
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:137:26  */
  /* ../neorv32/rtl/core/neorv32_cpu_regfile.vhd:134:20  */
endmodule

module neorv32_cpu_control_32_2_0_4_0_40_8cd82fcc1d144656bad81224642c94d0248852b6
  (input  clk_i,
   input  rstn_i,
   input  [31:0] i_bus_rdata_i,
   input  i_bus_ack_i,
   input  i_bus_err_i,
   input  i_pmp_fault_i,
   input  alu_cp_done_i,
   input  alu_exc_i,
   input  bus_d_wait_i,
   input  [1:0] cmp_i,
   input  [31:0] alu_add_i,
   input  [31:0] rs1_i,
   input  [4:0] fpu_flags_i,
   input  db_halt_req_i,
   input  msw_irq_i,
   input  mext_irq_i,
   input  mtime_irq_i,
   input  [15:0] firq_i,
   input  [31:0] mar_i,
   input  ma_load_i,
   input  ma_store_i,
   input  be_load_i,
   input  be_store_i,
   output ctrl_o_rf_wb_en,
   output [4:0] ctrl_o_rf_rs1,
   output [4:0] ctrl_o_rf_rs2,
   output [4:0] ctrl_o_rf_rs3,
   output [4:0] ctrl_o_rf_rd,
   output [1:0] ctrl_o_rf_mux,
   output ctrl_o_rf_zero_we,
   output [2:0] ctrl_o_alu_op,
   output ctrl_o_alu_opa_mux,
   output ctrl_o_alu_opb_mux,
   output ctrl_o_alu_unsigned,
   output [2:0] ctrl_o_alu_frm,
   output [5:0] ctrl_o_alu_cp_trig,
   output ctrl_o_bus_req,
   output ctrl_o_bus_mo_we,
   output ctrl_o_bus_fence,
   output ctrl_o_bus_fencei,
   output ctrl_o_bus_priv,
   output [2:0] ctrl_o_ir_funct3,
   output [11:0] ctrl_o_ir_funct12,
   output [6:0] ctrl_o_ir_opcode,
   output ctrl_o_cpu_priv,
   output ctrl_o_cpu_sleep,
   output ctrl_o_cpu_trap,
   output ctrl_o_cpu_debug,
   output [31:0] i_bus_addr_o,
   output i_bus_re_o,
   output [31:0] imm_o,
   output [31:0] curr_pc_o,
   output [31:0] next_pc_o,
   output [31:0] csr_rdata_o,
   output [543:0] pmp_addr_o,
   output [127:0] pmp_ctrl_o);
  wire n2756_o;
  wire [4:0] n2757_o;
  wire [4:0] n2758_o;
  wire [4:0] n2759_o;
  wire [4:0] n2760_o;
  wire [1:0] n2761_o;
  wire n2762_o;
  wire [2:0] n2763_o;
  wire n2764_o;
  wire n2765_o;
  wire n2766_o;
  wire [2:0] n2767_o;
  wire [5:0] n2768_o;
  wire n2769_o;
  wire n2770_o;
  wire n2771_o;
  wire n2772_o;
  wire n2773_o;
  wire [2:0] n2774_o;
  wire [11:0] n2775_o;
  wire [6:0] n2776_o;
  wire n2777_o;
  wire n2778_o;
  wire n2779_o;
  wire n2780_o;
  wire [41:0] fetch_engine;
  wire [79:0] ipb;
  wire [89:0] issue_engine;
  wire [7:0] decode_aux;
  wire [218:0] execute_engine;
  wire [101:0] trap_ctrl;
  wire [69:0] ctrl_nxt;
  wire [69:0] ctrl;
  wire [497:0] csr;
  wire [3231:0] cnt;
  wire [1023:0] cnt_lo_rd;
  wire [1023:0] cnt_hi_rd;
  wire [14:0] cnt_event;
  wire [8:0] debug_ctrl;
  wire illegal_cmd;
  wire csr_reg_valid;
  wire csr_rw_valid;
  wire csr_priv_valid;
  wire hw_trigger_fire;
  wire [6:0] imm_opcode;
  wire [11:0] csr_raddr;
  wire n2790_o;
  wire [1:0] n2798_o;
  wire [1:0] n2799_o;
  wire n2801_o;
  wire n2803_o;
  wire n2804_o;
  wire n2805_o;
  wire n2806_o;
  wire [1:0] n2807_o;
  wire [29:0] n2808_o;
  wire [31:0] n2810_o;
  wire n2811_o;
  wire n2814_o;
  wire [1:0] n2815_o;
  wire n2817_o;
  wire [1:0] n2819_o;
  wire [1:0] n2820_o;
  wire n2822_o;
  wire n2823_o;
  wire [31:0] n2824_o;
  wire [31:0] n2826_o;
  wire n2829_o;
  wire n2830_o;
  wire n2831_o;
  wire [4:0] n2833_o;
  wire n2835_o;
  wire n2836_o;
  wire n2837_o;
  wire [4:0] n2838_o;
  wire n2840_o;
  wire n2841_o;
  wire [4:0] n2842_o;
  wire n2844_o;
  wire n2845_o;
  wire [1:0] n2848_o;
  wire [1:0] n2849_o;
  wire [32:0] n2850_o;
  wire [1:0] n2851_o;
  wire [1:0] n2852_o;
  wire [32:0] n2853_o;
  wire [32:0] n2854_o;
  wire n2855_o;
  wire n2856_o;
  wire n2858_o;
  wire n2859_o;
  wire n2860_o;
  wire n2861_o;
  wire [1:0] n2864_o;
  wire n2866_o;
  wire [3:0] n2868_o;
  reg [1:0] n2869_o;
  wire n2870_o;
  wire n2871_o;
  reg n2872_o;
  wire [31:0] n2873_o;
  wire [31:0] n2874_o;
  reg [31:0] n2875_o;
  wire n2876_o;
  reg n2877_o;
  wire [37:0] n2878_o;
  wire [37:0] n2883_o;
  wire [29:0] n2887_o;
  wire [31:0] n2889_o;
  wire [1:0] n2891_o;
  wire n2893_o;
  wire [1:0] n2894_o;
  wire n2896_o;
  wire n2897_o;
  wire n2898_o;
  wire n2903_o;
  wire n2906_o;
  wire n2907_o;
  wire n2909_o;
  wire n2910_o;
  wire n2911_o;
  wire [1:0] n2912_o;
  wire [15:0] n2913_o;
  wire [17:0] n2914_o;
  wire n2915_o;
  wire n2916_o;
  wire n2917_o;
  wire [1:0] n2918_o;
  wire [15:0] n2919_o;
  wire [17:0] n2920_o;
  wire [1:0] n2922_o;
  wire n2924_o;
  wire n2925_o;
  wire n2926_o;
  wire n2927_o;
  wire n2928_o;
  wire n2930_o;
  wire n2931_o;
  wire n2932_o;
  wire [1:0] n2935_o;
  wire n2937_o;
  wire n2938_o;
  wire n2939_o;
  wire n2940_o;
  wire n2942_o;
  wire [17:0] n2944_o;
  wire n2945_o;
  wire prefetch_buffer_n1_prefetch_buffer_inst_n2946;
  wire n2947_o;
  wire [17:0] prefetch_buffer_n1_prefetch_buffer_inst_n2948;
  wire prefetch_buffer_n1_prefetch_buffer_inst_n2949;
  wire prefetch_buffer_n1_prefetch_buffer_inst_half_o;
  wire prefetch_buffer_n1_prefetch_buffer_inst_free_o;
  wire [17:0] prefetch_buffer_n1_prefetch_buffer_inst_rdata_o;
  wire prefetch_buffer_n1_prefetch_buffer_inst_avail_o;
  wire n2957_o;
  wire [17:0] n2959_o;
  wire n2960_o;
  wire prefetch_buffer_n2_prefetch_buffer_inst_n2961;
  wire n2962_o;
  wire [17:0] prefetch_buffer_n2_prefetch_buffer_inst_n2963;
  wire prefetch_buffer_n2_prefetch_buffer_inst_n2964;
  wire prefetch_buffer_n2_prefetch_buffer_inst_half_o;
  wire prefetch_buffer_n2_prefetch_buffer_inst_free_o;
  wire [17:0] prefetch_buffer_n2_prefetch_buffer_inst_rdata_o;
  wire prefetch_buffer_n2_prefetch_buffer_inst_avail_o;
  wire n2974_o;
  wire n2975_o;
  wire [3:0] n2976_o;
  wire n2978_o;
  wire n2979_o;
  wire n2980_o;
  wire n2981_o;
  wire n2982_o;
  wire n2983_o;
  wire n2984_o;
  wire n2985_o;
  wire n2986_o;
  wire n2987_o;
  localparam [1:0] n2994_o = 2'b00;
  wire n2995_o;
  wire n2996_o;
  wire [1:0] n2997_o;
  wire n2999_o;
  wire n3000_o;
  wire n3001_o;
  wire n3002_o;
  wire [1:0] n3003_o;
  wire [2:0] n3004_o;
  wire [3:0] n3006_o;
  wire [31:0] n3007_o;
  wire [35:0] n3008_o;
  wire n3009_o;
  wire n3010_o;
  wire n3011_o;
  wire n3012_o;
  wire n3013_o;
  wire n3014_o;
  wire [1:0] n3015_o;
  wire [1:0] n3016_o;
  wire [1:0] n3017_o;
  wire [1:0] n3018_o;
  wire [2:0] n3020_o;
  wire [3:0] n3022_o;
  wire [15:0] n3023_o;
  wire [15:0] n3024_o;
  wire [31:0] n3025_o;
  wire [35:0] n3026_o;
  wire [37:0] n3027_o;
  wire [36:0] n3028_o;
  wire n3029_o;
  wire [36:0] n3030_o;
  wire [36:0] n3031_o;
  wire n3032_o;
  wire n3033_o;
  wire n3034_o;
  wire [1:0] n3035_o;
  wire n3037_o;
  wire n3038_o;
  wire n3039_o;
  wire n3040_o;
  wire [1:0] n3041_o;
  wire [2:0] n3042_o;
  wire [3:0] n3044_o;
  wire [31:0] n3045_o;
  wire [35:0] n3046_o;
  wire n3047_o;
  wire n3048_o;
  wire n3049_o;
  wire n3050_o;
  wire n3051_o;
  wire n3052_o;
  wire [1:0] n3053_o;
  wire [1:0] n3054_o;
  wire [1:0] n3055_o;
  wire [1:0] n3056_o;
  wire [2:0] n3058_o;
  wire [3:0] n3060_o;
  wire [15:0] n3061_o;
  wire [15:0] n3062_o;
  wire [31:0] n3063_o;
  wire [35:0] n3064_o;
  wire [37:0] n3065_o;
  wire n3066_o;
  wire [35:0] n3067_o;
  wire [35:0] n3068_o;
  wire n3069_o;
  wire n3070_o;
  wire n3071_o;
  wire n3072_o;
  wire n3073_o;
  wire [37:0] n3074_o;
  wire [37:0] n3075_o;
  wire n3076_o;
  wire n3077_o;
  wire [37:0] n3078_o;
  wire n3081_o;
  wire [3:0] n3082_o;
  wire n3084_o;
  wire n3085_o;
  wire n3086_o;
  wire n3089_o;
  wire [3:0] n3090_o;
  wire n3092_o;
  wire n3093_o;
  wire n3094_o;
  wire [15:0] n3096_o;
  wire neorv32_cpu_decompressor_inst_true_neorv32_cpu_decompressor_inst_n3097;
  wire [31:0] neorv32_cpu_decompressor_inst_true_neorv32_cpu_decompressor_inst_n3098;
  wire neorv32_cpu_decompressor_inst_true_neorv32_cpu_decompressor_inst_ci_illegal_o;
  wire [31:0] neorv32_cpu_decompressor_inst_true_neorv32_cpu_decompressor_inst_ci_instr32_o;
  wire [15:0] n3103_o;
  wire n3104_o;
  wire n3105_o;
  wire [15:0] n3106_o;
  wire [15:0] n3107_o;
  wire n3110_o;
  wire n3111_o;
  wire n3112_o;
  wire n3113_o;
  wire n3114_o;
  wire n3115_o;
  wire n3116_o;
  wire n3117_o;
  wire n3118_o;
  wire n3119_o;
  wire n3120_o;
  wire n3121_o;
  wire n3122_o;
  wire n3123_o;
  wire n3124_o;
  wire n3125_o;
  wire n3126_o;
  wire n3127_o;
  wire n3128_o;
  wire n3129_o;
  wire n3130_o;
  wire [3:0] n3131_o;
  wire [3:0] n3132_o;
  wire [3:0] n3133_o;
  wire [3:0] n3134_o;
  wire [3:0] n3135_o;
  wire [15:0] n3136_o;
  wire [4:0] n3137_o;
  wire [20:0] n3138_o;
  wire [5:0] n3139_o;
  wire [4:0] n3140_o;
  wire n3142_o;
  wire n3143_o;
  wire n3144_o;
  wire n3145_o;
  wire n3146_o;
  wire n3147_o;
  wire n3148_o;
  wire n3149_o;
  wire n3150_o;
  wire n3151_o;
  wire n3152_o;
  wire n3153_o;
  wire n3154_o;
  wire n3155_o;
  wire n3156_o;
  wire n3157_o;
  wire n3158_o;
  wire n3159_o;
  wire n3160_o;
  wire n3161_o;
  wire n3162_o;
  wire [3:0] n3163_o;
  wire [3:0] n3164_o;
  wire [3:0] n3165_o;
  wire [3:0] n3166_o;
  wire [3:0] n3167_o;
  wire [15:0] n3168_o;
  wire [19:0] n3169_o;
  wire n3170_o;
  wire [5:0] n3171_o;
  wire [3:0] n3172_o;
  wire n3175_o;
  wire [19:0] n3176_o;
  localparam [11:0] n3177_o = 12'b000000000000;
  wire n3179_o;
  wire n3181_o;
  wire n3182_o;
  wire n3183_o;
  wire n3184_o;
  wire n3185_o;
  wire n3186_o;
  wire n3187_o;
  wire n3188_o;
  wire n3189_o;
  wire n3190_o;
  wire n3191_o;
  wire n3192_o;
  wire n3193_o;
  wire n3194_o;
  wire [3:0] n3195_o;
  wire [3:0] n3196_o;
  wire [3:0] n3197_o;
  wire [11:0] n3198_o;
  wire [7:0] n3199_o;
  wire n3200_o;
  wire [9:0] n3201_o;
  wire n3204_o;
  wire n3205_o;
  wire n3206_o;
  wire n3207_o;
  wire n3208_o;
  wire n3209_o;
  wire n3210_o;
  wire n3211_o;
  wire n3212_o;
  wire n3213_o;
  wire n3214_o;
  wire n3215_o;
  wire n3216_o;
  wire n3217_o;
  wire n3218_o;
  wire n3219_o;
  wire n3220_o;
  wire n3221_o;
  wire n3222_o;
  wire n3223_o;
  wire n3224_o;
  wire n3225_o;
  wire [3:0] n3226_o;
  wire [3:0] n3227_o;
  wire [3:0] n3228_o;
  wire [3:0] n3229_o;
  wire [3:0] n3230_o;
  wire [15:0] n3231_o;
  wire [4:0] n3232_o;
  wire [20:0] n3233_o;
  wire [9:0] n3234_o;
  wire n3235_o;
  wire [3:0] n3236_o;
  wire n3237_o;
  wire n3238_o;
  reg n3239_o;
  wire [3:0] n3240_o;
  wire [3:0] n3241_o;
  wire [3:0] n3242_o;
  wire [3:0] n3243_o;
  reg [3:0] n3244_o;
  wire [5:0] n3245_o;
  wire [5:0] n3246_o;
  wire [5:0] n3247_o;
  reg [5:0] n3248_o;
  wire n3249_o;
  wire n3250_o;
  wire n3251_o;
  reg n3252_o;
  wire [7:0] n3253_o;
  wire [7:0] n3254_o;
  wire [7:0] n3255_o;
  wire [7:0] n3256_o;
  reg [7:0] n3257_o;
  wire [11:0] n3258_o;
  wire [11:0] n3259_o;
  wire [11:0] n3260_o;
  wire [11:0] n3261_o;
  reg [11:0] n3262_o;
  wire [31:0] n3263_o;
  wire [4:0] n3266_o;
  wire [6:0] n3268_o;
  wire n3270_o;
  wire n3271_o;
  wire n3272_o;
  wire n3273_o;
  wire n3274_o;
  wire n3275_o;
  wire n3276_o;
  wire n3277_o;
  wire n3278_o;
  wire n3281_o;
  wire [3:0] n3294_o;
  wire [3:0] n3295_o;
  wire [3:0] n3296_o;
  wire n3297_o;
  wire [31:0] n3298_o;
  wire n3299_o;
  wire n3300_o;
  wire n3301_o;
  wire [3:0] n3302_o;
  wire n3304_o;
  wire [31:0] n3305_o;
  wire [31:0] n3306_o;
  wire [31:0] n3307_o;
  wire n3308_o;
  wire n3309_o;
  wire n3310_o;
  wire [30:0] n3311_o;
  wire [31:0] n3313_o;
  wire [30:0] n3314_o;
  wire [31:0] n3316_o;
  wire [31:0] n3317_o;
  wire [3:0] n3320_o;
  wire [29:0] n3323_o;
  wire [31:0] n3325_o;
  wire n3327_o;
  wire [30:0] n3329_o;
  wire [31:0] n3331_o;
  wire n3333_o;
  wire [31:0] n3334_o;
  wire [31:0] n3335_o;
  wire [31:0] n3336_o;
  wire n3338_o;
  wire [2:0] n3339_o;
  wire [31:0] n3340_o;
  reg [31:0] n3341_o;
  wire [39:0] n3342_o;
  wire [32:0] n3343_o;
  wire [39:0] n3361_o;
  wire [32:0] n3362_o;
  wire n3376_o;
  wire n3377_o;
  wire n3379_o;
  wire [3:0] n3380_o;
  wire [30:0] n3382_o;
  wire [31:0] n3384_o;
  wire [30:0] n3385_o;
  wire [31:0] n3387_o;
  wire n3389_o;
  wire n3390_o;
  wire n3391_o;
  wire n3392_o;
  wire [4:0] n3393_o;
  wire [4:0] n3394_o;
  wire [4:0] n3395_o;
  wire [4:0] n3396_o;
  wire [1:0] n3397_o;
  wire n3398_o;
  wire [2:0] n3399_o;
  wire n3400_o;
  wire n3401_o;
  wire n3402_o;
  wire [2:0] n3403_o;
  wire [5:0] n3404_o;
  wire n3405_o;
  wire n3406_o;
  wire n3407_o;
  wire n3408_o;
  wire n3409_o;
  wire n3410_o;
  wire n3411_o;
  wire n3412_o;
  wire [2:0] n3413_o;
  wire [11:0] n3414_o;
  wire [6:0] n3415_o;
  wire n3416_o;
  wire n3417_o;
  wire n3418_o;
  wire n3419_o;
  wire [6:0] n3430_o;
  wire n3432_o;
  wire n3433_o;
  wire n3434_o;
  wire n3436_o;
  wire n3438_o;
  wire n3439_o;
  wire n3441_o;
  wire n3443_o;
  wire [1:0] n3444_o;
  wire [1:0] n3445_o;
  wire [1:0] n3446_o;
  wire [4:0] n3447_o;
  wire n3449_o;
  wire n3451_o;
  wire [4:0] n3452_o;
  wire n3454_o;
  wire n3456_o;
  wire [11:0] n3458_o;
  wire [3:0] n3460_o;
  wire [31:0] n3461_o;
  wire n3462_o;
  wire n3464_o;
  wire n3465_o;
  localparam [69:0] n3479_o = 70'b0000000000000000000000000000000000000000000000000000000000000000000000;
  wire n3483_o;
  wire n3485_o;
  wire n3486_o;
  wire n3487_o;
  wire n3488_o;
  wire [3:0] n3491_o;
  wire n3493_o;
  wire n3494_o;
  wire n3495_o;
  wire n3496_o;
  wire n3497_o;
  wire n3498_o;
  wire n3499_o;
  wire [31:0] n3500_o;
  wire n3502_o;
  wire n3505_o;
  wire n3506_o;
  wire n3507_o;
  wire n3508_o;
  wire n3509_o;
  wire n3510_o;
  wire n3511_o;
  wire n3514_o;
  wire n3515_o;
  wire n3516_o;
  wire [3:0] n3519_o;
  wire [3:0] n3520_o;
  wire [31:0] n3521_o;
  wire n3522_o;
  wire [1:0] n3523_o;
  wire [1:0] n3524_o;
  wire [1:0] n3525_o;
  wire n3527_o;
  wire n3528_o;
  wire [3:0] n3531_o;
  wire n3532_o;
  wire n3534_o;
  wire n3538_o;
  wire n3545_o;
  wire [6:0] n3546_o;
  wire n3547_o;
  wire n3548_o;
  wire n3550_o;
  wire n3551_o;
  wire [2:0] n3552_o;
  wire n3553_o;
  wire n3554_o;
  wire n3555_o;
  wire [2:0] n3557_o;
  wire n3559_o;
  wire n3562_o;
  wire n3564_o;
  wire n3565_o;
  wire n3568_o;
  wire n3571_o;
  wire [3:0] n3573_o;
  reg [2:0] n3574_o;
  wire n3575_o;
  wire n3577_o;
  wire n3578_o;
  wire n3579_o;
  wire n3580_o;
  wire n3581_o;
  wire n3583_o;
  wire [2:0] n3586_o;
  wire n3588_o;
  wire [2:0] n3589_o;
  wire n3591_o;
  wire n3592_o;
  wire [3:0] n3597_o;
  wire n3598_o;
  wire n3599_o;
  wire n3600_o;
  wire n3601_o;
  wire [3:0] n3602_o;
  wire n3603_o;
  wire n3604_o;
  wire n3605_o;
  wire n3606_o;
  wire n3607_o;
  wire n3608_o;
  wire n3610_o;
  wire n3612_o;
  wire n3613_o;
  wire n3616_o;
  wire [2:0] n3618_o;
  wire n3622_o;
  wire n3624_o;
  wire n3625_o;
  wire n3630_o;
  wire n3632_o;
  wire n3633_o;
  wire [1:0] n3635_o;
  wire n3637_o;
  wire n3640_o;
  wire n3643_o;
  wire n3645_o;
  wire n3646_o;
  wire n3648_o;
  wire n3649_o;
  wire [2:0] n3650_o;
  wire n3652_o;
  wire n3654_o;
  wire n3655_o;
  wire n3661_o;
  wire n3664_o;
  wire n3667_o;
  wire n3669_o;
  wire n3670_o;
  wire n3672_o;
  wire n3673_o;
  wire n3675_o;
  wire n3676_o;
  wire n3680_o;
  wire [7:0] n3682_o;
  reg [3:0] n3683_o;
  wire n3684_o;
  reg n3685_o;
  reg [2:0] n3686_o;
  wire n3687_o;
  reg n3688_o;
  wire n3689_o;
  reg n3690_o;
  wire n3691_o;
  reg n3692_o;
  wire n3693_o;
  reg n3694_o;
  wire n3695_o;
  reg n3696_o;
  wire n3697_o;
  reg n3698_o;
  reg n3699_o;
  wire n3701_o;
  wire n3703_o;
  wire n3704_o;
  wire [3:0] n3707_o;
  wire n3708_o;
  wire n3709_o;
  wire n3711_o;
  wire n3715_o;
  wire n3716_o;
  wire n3717_o;
  wire n3721_o;
  wire [3:0] n3722_o;
  wire n3723_o;
  wire n3725_o;
  wire n3726_o;
  wire n3728_o;
  wire n3734_o;
  wire n3735_o;
  wire n3736_o;
  wire n3738_o;
  wire n3739_o;
  wire n3742_o;
  wire n3744_o;
  wire n3745_o;
  wire n3746_o;
  wire n3747_o;
  wire n3748_o;
  wire n3749_o;
  wire n3750_o;
  wire n3751_o;
  wire n3752_o;
  wire n3754_o;
  wire n3755_o;
  wire n3756_o;
  wire n3758_o;
  wire n3759_o;
  wire [3:0] n3761_o;
  wire n3763_o;
  wire [3:0] n3764_o;
  wire n3765_o;
  wire n3766_o;
  wire n3768_o;
  wire [2:0] n3769_o;
  wire n3771_o;
  wire n3772_o;
  wire n3773_o;
  wire n3774_o;
  wire [11:0] n3776_o;
  wire n3779_o;
  wire n3782_o;
  wire n3785_o;
  wire n3789_o;
  wire [3:0] n3791_o;
  reg [3:0] n3792_o;
  reg n3793_o;
  reg n3794_o;
  reg n3795_o;
  reg n3796_o;
  wire [2:0] n3798_o;
  wire n3800_o;
  wire [2:0] n3801_o;
  wire n3803_o;
  wire n3804_o;
  wire n3805_o;
  wire n3806_o;
  wire n3807_o;
  wire n3809_o;
  wire [3:0] n3811_o;
  wire n3812_o;
  wire [1:0] n3813_o;
  wire [1:0] n3814_o;
  wire [1:0] n3815_o;
  wire n3816_o;
  wire n3817_o;
  wire n3818_o;
  wire n3819_o;
  wire n3821_o;
  wire [10:0] n3823_o;
  reg n3824_o;
  reg [3:0] n3825_o;
  reg [31:0] n3826_o;
  reg n3827_o;
  reg n3828_o;
  reg n3829_o;
  reg n3830_o;
  reg n3831_o;
  reg n3832_o;
  reg n3833_o;
  reg n3834_o;
  wire [1:0] n3835_o;
  reg [1:0] n3836_o;
  wire [1:0] n3837_o;
  reg [1:0] n3838_o;
  wire n3839_o;
  reg n3840_o;
  reg [1:0] n3841_o;
  reg n3842_o;
  reg [2:0] n3843_o;
  wire n3844_o;
  reg n3845_o;
  wire n3846_o;
  reg n3847_o;
  wire n3848_o;
  reg n3849_o;
  wire n3850_o;
  reg n3851_o;
  wire n3852_o;
  reg n3853_o;
  wire n3854_o;
  reg n3855_o;
  wire n3856_o;
  reg n3857_o;
  wire [19:0] n3858_o;
  wire [2:0] n3861_o;
  wire [3:0] n3864_o;
  wire [27:0] n3866_o;
  reg n3867_o;
  reg n3868_o;
  reg n3869_o;
  wire [11:0] n3872_o;
  wire n3875_o;
  wire n3877_o;
  wire n3878_o;
  wire n3880_o;
  wire n3881_o;
  wire n3883_o;
  wire n3885_o;
  wire n3886_o;
  wire n3888_o;
  wire n3889_o;
  wire n3891_o;
  wire n3892_o;
  wire n3894_o;
  wire n3895_o;
  wire n3897_o;
  wire n3898_o;
  wire n3900_o;
  wire n3901_o;
  wire n3903_o;
  wire n3904_o;
  wire n3906_o;
  wire n3907_o;
  wire n3909_o;
  wire n3910_o;
  wire n3912_o;
  wire n3913_o;
  wire n3915_o;
  wire n3916_o;
  wire n3918_o;
  wire n3919_o;
  wire n3921_o;
  wire n3922_o;
  wire n3924_o;
  wire n3925_o;
  wire n3927_o;
  wire n3928_o;
  wire n3930_o;
  wire n3931_o;
  wire n3933_o;
  wire n3934_o;
  wire n3936_o;
  wire n3937_o;
  wire n3939_o;
  wire n3940_o;
  wire n3943_o;
  wire n3945_o;
  wire n3946_o;
  wire n3948_o;
  wire n3949_o;
  wire n3951_o;
  wire n3952_o;
  wire n3954_o;
  wire n3955_o;
  wire n3957_o;
  wire n3958_o;
  wire n3960_o;
  wire n3961_o;
  wire n3963_o;
  wire n3964_o;
  wire n3966_o;
  wire n3967_o;
  wire n3969_o;
  wire n3970_o;
  wire n3972_o;
  wire n3973_o;
  wire n3975_o;
  wire n3976_o;
  wire n3978_o;
  wire n3979_o;
  wire n3981_o;
  wire n3982_o;
  wire n3984_o;
  wire n3985_o;
  wire n3987_o;
  wire n3988_o;
  wire n3990_o;
  wire n3991_o;
  wire n3993_o;
  wire n3994_o;
  wire n3996_o;
  wire n3997_o;
  wire n3999_o;
  wire n4000_o;
  wire n4003_o;
  wire n4005_o;
  wire n4006_o;
  wire n4008_o;
  wire n4009_o;
  wire n4011_o;
  wire n4012_o;
  wire n4014_o;
  wire n4015_o;
  wire n4017_o;
  wire n4018_o;
  wire n4020_o;
  wire n4021_o;
  wire n4023_o;
  wire n4024_o;
  wire n4026_o;
  wire n4027_o;
  wire n4029_o;
  wire n4030_o;
  wire n4032_o;
  wire n4033_o;
  wire n4035_o;
  wire n4036_o;
  wire n4038_o;
  wire n4039_o;
  wire n4041_o;
  wire n4042_o;
  wire n4044_o;
  wire n4045_o;
  wire n4047_o;
  wire n4048_o;
  wire n4050_o;
  wire n4051_o;
  wire n4053_o;
  wire n4054_o;
  wire n4056_o;
  wire n4057_o;
  wire n4059_o;
  wire n4060_o;
  wire n4062_o;
  wire n4063_o;
  wire n4065_o;
  wire n4066_o;
  wire n4068_o;
  wire n4069_o;
  wire n4071_o;
  wire n4072_o;
  wire n4074_o;
  wire n4075_o;
  wire n4077_o;
  wire n4078_o;
  wire n4080_o;
  wire n4081_o;
  wire n4083_o;
  wire n4084_o;
  wire n4086_o;
  wire n4087_o;
  wire n4089_o;
  wire n4090_o;
  wire n4092_o;
  wire n4093_o;
  wire n4095_o;
  wire n4096_o;
  wire n4098_o;
  wire n4099_o;
  wire n4101_o;
  wire n4102_o;
  wire n4104_o;
  wire n4105_o;
  wire n4107_o;
  wire n4108_o;
  wire n4110_o;
  wire n4111_o;
  wire n4113_o;
  wire n4114_o;
  wire n4116_o;
  wire n4117_o;
  wire n4119_o;
  wire n4120_o;
  wire n4122_o;
  wire n4123_o;
  wire n4125_o;
  wire n4126_o;
  wire n4128_o;
  wire n4129_o;
  wire n4131_o;
  wire n4132_o;
  wire n4134_o;
  wire n4135_o;
  wire n4137_o;
  wire n4138_o;
  wire n4140_o;
  wire n4141_o;
  wire n4143_o;
  wire n4144_o;
  wire n4146_o;
  wire n4147_o;
  wire n4149_o;
  wire n4150_o;
  wire n4152_o;
  wire n4153_o;
  wire n4155_o;
  wire n4156_o;
  wire n4158_o;
  wire n4159_o;
  wire n4161_o;
  wire n4162_o;
  wire n4164_o;
  wire n4165_o;
  wire n4167_o;
  wire n4168_o;
  wire n4170_o;
  wire n4171_o;
  wire n4173_o;
  wire n4174_o;
  wire n4176_o;
  wire n4177_o;
  wire n4179_o;
  wire n4180_o;
  wire n4182_o;
  wire n4183_o;
  wire n4185_o;
  wire n4186_o;
  wire n4188_o;
  wire n4189_o;
  wire n4191_o;
  wire n4192_o;
  wire n4194_o;
  wire n4195_o;
  wire n4197_o;
  wire n4198_o;
  wire n4200_o;
  wire n4201_o;
  wire n4203_o;
  wire n4204_o;
  wire n4206_o;
  wire n4207_o;
  wire n4209_o;
  wire n4210_o;
  wire n4212_o;
  wire n4213_o;
  wire n4215_o;
  wire n4216_o;
  wire n4218_o;
  wire n4219_o;
  wire n4221_o;
  wire n4222_o;
  wire n4224_o;
  wire n4225_o;
  wire n4227_o;
  wire n4228_o;
  wire n4230_o;
  wire n4231_o;
  wire n4233_o;
  wire n4234_o;
  wire n4236_o;
  wire n4237_o;
  wire n4239_o;
  wire n4240_o;
  wire n4242_o;
  wire n4243_o;
  wire n4245_o;
  wire n4246_o;
  wire n4248_o;
  wire n4249_o;
  wire n4251_o;
  wire n4252_o;
  wire n4254_o;
  wire n4255_o;
  wire n4257_o;
  wire n4258_o;
  wire n4260_o;
  wire n4261_o;
  wire n4263_o;
  wire n4264_o;
  wire n4266_o;
  wire n4267_o;
  wire n4269_o;
  wire n4270_o;
  wire n4272_o;
  wire n4273_o;
  wire n4275_o;
  wire n4276_o;
  wire n4278_o;
  wire n4279_o;
  wire n4281_o;
  wire n4282_o;
  wire n4284_o;
  wire n4285_o;
  wire n4287_o;
  wire n4288_o;
  wire n4290_o;
  wire n4291_o;
  wire n4293_o;
  wire n4294_o;
  wire n4296_o;
  wire n4297_o;
  wire n4299_o;
  wire n4300_o;
  wire n4302_o;
  wire n4303_o;
  wire n4305_o;
  wire n4306_o;
  wire n4308_o;
  wire n4309_o;
  wire n4311_o;
  wire n4312_o;
  wire n4314_o;
  wire n4315_o;
  wire n4317_o;
  wire n4318_o;
  wire n4320_o;
  wire n4321_o;
  wire n4323_o;
  wire n4324_o;
  wire n4326_o;
  wire n4327_o;
  wire n4329_o;
  wire n4330_o;
  wire n4332_o;
  wire n4333_o;
  wire n4335_o;
  wire n4336_o;
  wire n4338_o;
  wire n4339_o;
  wire n4341_o;
  wire n4342_o;
  wire n4344_o;
  wire n4345_o;
  wire n4347_o;
  wire n4348_o;
  wire n4350_o;
  wire n4351_o;
  wire n4353_o;
  wire n4354_o;
  wire n4356_o;
  wire n4357_o;
  wire n4359_o;
  wire n4360_o;
  wire n4362_o;
  wire n4363_o;
  wire n4365_o;
  wire n4366_o;
  wire n4368_o;
  wire n4369_o;
  wire n4371_o;
  wire n4372_o;
  wire n4374_o;
  wire n4375_o;
  wire n4377_o;
  wire n4378_o;
  wire n4380_o;
  wire n4381_o;
  wire n4383_o;
  wire n4384_o;
  wire n4386_o;
  wire n4387_o;
  wire n4389_o;
  wire n4390_o;
  wire n4392_o;
  wire n4393_o;
  wire n4395_o;
  wire n4396_o;
  wire n4398_o;
  wire n4399_o;
  wire n4401_o;
  wire n4402_o;
  wire n4404_o;
  wire n4405_o;
  wire n4407_o;
  wire n4408_o;
  wire n4410_o;
  wire n4411_o;
  wire n4413_o;
  wire n4414_o;
  wire n4416_o;
  wire n4417_o;
  wire n4419_o;
  wire n4420_o;
  wire n4422_o;
  wire n4423_o;
  wire n4425_o;
  wire n4426_o;
  wire n4428_o;
  wire n4429_o;
  wire n4431_o;
  wire n4432_o;
  wire n4434_o;
  wire n4435_o;
  wire n4438_o;
  wire n4440_o;
  wire n4441_o;
  wire n4443_o;
  wire n4444_o;
  wire n4446_o;
  wire n4447_o;
  wire n4449_o;
  wire n4450_o;
  wire n4452_o;
  wire n4453_o;
  wire n4455_o;
  wire n4456_o;
  wire n4458_o;
  wire n4459_o;
  wire n4461_o;
  wire n4462_o;
  wire n4464_o;
  wire n4465_o;
  wire n4468_o;
  wire n4470_o;
  wire n4471_o;
  wire n4473_o;
  wire n4474_o;
  wire n4477_o;
  wire n4479_o;
  wire n4480_o;
  wire n4482_o;
  wire n4483_o;
  wire n4485_o;
  wire n4486_o;
  wire n4488_o;
  wire n4489_o;
  wire n4491_o;
  wire n4492_o;
  wire n4494_o;
  wire n4495_o;
  wire n4497_o;
  wire n4498_o;
  wire [6:0] n4499_o;
  reg n4508_o;
  wire [1:0] n4512_o;
  wire n4514_o;
  wire [2:0] n4515_o;
  wire n4517_o;
  wire [2:0] n4518_o;
  wire n4520_o;
  wire n4521_o;
  wire n4522_o;
  wire n4523_o;
  wire n4524_o;
  wire n4525_o;
  wire n4528_o;
  wire [1:0] n4547_o;
  wire n4549_o;
  wire n4550_o;
  wire n4551_o;
  wire n4552_o;
  wire n4555_o;
  wire [6:0] n4558_o;
  wire n4560_o;
  wire n4562_o;
  wire n4563_o;
  wire n4565_o;
  wire n4566_o;
  wire [2:0] n4567_o;
  wire n4569_o;
  reg n4572_o;
  wire n4574_o;
  wire [2:0] n4575_o;
  wire n4577_o;
  wire n4579_o;
  wire n4580_o;
  wire n4582_o;
  wire n4583_o;
  wire n4585_o;
  wire n4586_o;
  wire n4588_o;
  wire n4589_o;
  wire n4591_o;
  wire n4592_o;
  reg n4595_o;
  wire n4597_o;
  wire [2:0] n4598_o;
  wire n4600_o;
  wire n4602_o;
  wire n4603_o;
  wire n4605_o;
  wire n4606_o;
  wire n4608_o;
  wire n4609_o;
  wire n4611_o;
  wire n4612_o;
  reg n4615_o;
  wire n4617_o;
  wire [2:0] n4618_o;
  wire n4620_o;
  wire n4622_o;
  wire n4623_o;
  wire n4625_o;
  wire n4626_o;
  reg n4629_o;
  wire n4631_o;
  wire [2:0] n4632_o;
  wire n4634_o;
  wire [2:0] n4635_o;
  wire n4637_o;
  wire n4638_o;
  wire [4:0] n4639_o;
  wire n4641_o;
  wire n4642_o;
  wire n4643_o;
  wire n4644_o;
  wire n4645_o;
  wire [2:0] n4646_o;
  wire n4648_o;
  wire [2:0] n4649_o;
  wire n4651_o;
  wire n4652_o;
  wire [2:0] n4653_o;
  wire n4655_o;
  wire n4656_o;
  wire [2:0] n4657_o;
  wire n4659_o;
  wire n4660_o;
  wire [2:0] n4661_o;
  wire n4663_o;
  wire n4664_o;
  wire [2:0] n4665_o;
  wire n4667_o;
  wire n4668_o;
  wire [6:0] n4669_o;
  wire n4671_o;
  wire n4672_o;
  wire n4673_o;
  wire n4674_o;
  wire n4676_o;
  wire n4677_o;
  wire n4678_o;
  wire n4680_o;
  wire n4681_o;
  wire n4683_o;
  wire n4685_o;
  wire n4688_o;
  wire n4690_o;
  wire [2:0] n4691_o;
  wire n4693_o;
  wire [2:0] n4694_o;
  wire n4696_o;
  wire n4697_o;
  wire [2:0] n4698_o;
  wire n4700_o;
  wire n4701_o;
  wire [2:0] n4702_o;
  wire n4704_o;
  wire n4705_o;
  wire [2:0] n4706_o;
  wire n4708_o;
  wire n4709_o;
  wire [2:0] n4710_o;
  wire n4712_o;
  wire n4713_o;
  wire [2:0] n4714_o;
  wire n4716_o;
  wire [6:0] n4717_o;
  wire n4719_o;
  wire n4720_o;
  wire n4721_o;
  wire [2:0] n4722_o;
  wire n4724_o;
  wire [4:0] n4725_o;
  wire n4727_o;
  wire n4728_o;
  wire n4729_o;
  wire n4730_o;
  wire n4731_o;
  wire n4732_o;
  wire n4734_o;
  wire n4737_o;
  wire n4739_o;
  wire [2:0] n4740_o;
  wire n4742_o;
  wire n4745_o;
  wire [1:0] n4746_o;
  reg n4750_o;
  wire n4752_o;
  wire [2:0] n4753_o;
  wire n4755_o;
  wire n4756_o;
  wire n4757_o;
  wire n4758_o;
  wire [11:0] n4759_o;
  wire n4761_o;
  wire n4763_o;
  wire n4764_o;
  wire n4765_o;
  wire n4766_o;
  wire n4768_o;
  wire n4769_o;
  wire n4770_o;
  wire n4771_o;
  wire n4772_o;
  wire n4774_o;
  wire n4775_o;
  wire n4776_o;
  wire n4778_o;
  wire [3:0] n4779_o;
  reg n4782_o;
  wire n4784_o;
  wire n4785_o;
  wire n4786_o;
  wire n4787_o;
  wire n4788_o;
  wire n4789_o;
  wire [2:0] n4790_o;
  wire n4792_o;
  wire n4793_o;
  wire n4796_o;
  wire n4797_o;
  wire n4799_o;
  wire n4801_o;
  wire n4802_o;
  wire n4804_o;
  wire n4806_o;
  wire n4809_o;
  wire n4811_o;
  wire n4812_o;
  wire n4814_o;
  wire n4815_o;
  wire n4817_o;
  wire n4818_o;
  wire [10:0] n4819_o;
  reg n4823_o;
  wire n4826_o;
  wire n4828_o;
  wire n4830_o;
  wire n4831_o;
  wire [3:0] n4832_o;
  wire n4834_o;
  wire [3:0] n4835_o;
  wire n4837_o;
  wire n4838_o;
  wire n4839_o;
  wire n4842_o;
  wire n4847_o;
  wire n4848_o;
  wire n4849_o;
  wire n4850_o;
  wire n4851_o;
  wire n4852_o;
  wire n4853_o;
  wire n4854_o;
  wire n4855_o;
  wire n4856_o;
  wire n4857_o;
  wire n4858_o;
  wire n4859_o;
  wire n4860_o;
  wire n4861_o;
  wire n4862_o;
  wire n4863_o;
  wire n4864_o;
  wire n4865_o;
  wire n4866_o;
  wire n4867_o;
  wire n4868_o;
  wire n4869_o;
  wire n4870_o;
  wire n4871_o;
  wire n4872_o;
  wire n4873_o;
  wire n4874_o;
  wire n4875_o;
  wire n4876_o;
  wire n4877_o;
  wire n4878_o;
  wire n4879_o;
  wire n4880_o;
  wire n4881_o;
  wire n4882_o;
  wire n4883_o;
  wire n4884_o;
  wire n4885_o;
  wire n4886_o;
  wire n4887_o;
  wire n4888_o;
  wire n4889_o;
  wire n4890_o;
  wire n4891_o;
  wire n4892_o;
  wire n4893_o;
  wire n4894_o;
  wire n4895_o;
  wire n4896_o;
  wire n4897_o;
  wire n4900_o;
  wire n4901_o;
  wire n4902_o;
  wire n4903_o;
  wire n4904_o;
  wire n4905_o;
  wire n4906_o;
  wire n4907_o;
  wire n4908_o;
  wire n4909_o;
  wire n4910_o;
  wire n4911_o;
  wire n4912_o;
  wire n4913_o;
  wire n4914_o;
  wire n4915_o;
  wire n4916_o;
  wire n4917_o;
  wire n4918_o;
  wire n4919_o;
  wire n4920_o;
  wire n4921_o;
  wire n4922_o;
  wire n4923_o;
  wire n4924_o;
  wire n4925_o;
  wire n4926_o;
  wire n4927_o;
  wire n4928_o;
  wire n4929_o;
  wire n4930_o;
  wire n4931_o;
  wire n4932_o;
  wire n4933_o;
  wire n4934_o;
  wire n4935_o;
  wire n4936_o;
  wire n4937_o;
  wire n4938_o;
  wire n4939_o;
  wire n4940_o;
  wire n4941_o;
  wire n4942_o;
  wire n4943_o;
  wire n4944_o;
  wire n4945_o;
  wire n4946_o;
  wire n4947_o;
  wire n4948_o;
  wire n4949_o;
  wire n4950_o;
  wire n4951_o;
  wire n4952_o;
  wire n4953_o;
  wire n4954_o;
  wire n4955_o;
  wire n4956_o;
  wire n4957_o;
  wire n4958_o;
  wire n4959_o;
  wire n4960_o;
  wire n4961_o;
  wire n4962_o;
  wire n4963_o;
  wire n4964_o;
  wire n4965_o;
  wire n4966_o;
  wire n4967_o;
  wire n4968_o;
  wire n4969_o;
  wire n4970_o;
  wire n4971_o;
  wire n4972_o;
  wire n4973_o;
  wire n4974_o;
  wire n4975_o;
  wire n4976_o;
  wire n4977_o;
  wire n4978_o;
  wire n4979_o;
  wire n4982_o;
  wire n4983_o;
  wire n4984_o;
  wire n4985_o;
  wire n4986_o;
  wire n4987_o;
  wire n4988_o;
  wire n4989_o;
  wire n4990_o;
  wire n4991_o;
  wire n4992_o;
  wire n4993_o;
  wire n4994_o;
  wire n4995_o;
  wire n4996_o;
  wire n4997_o;
  wire n4998_o;
  wire n4999_o;
  wire n5000_o;
  wire n5001_o;
  wire n5002_o;
  wire n5003_o;
  wire n5004_o;
  wire n5005_o;
  wire n5006_o;
  wire n5007_o;
  wire n5008_o;
  wire n5009_o;
  wire n5010_o;
  wire n5011_o;
  wire n5012_o;
  wire n5013_o;
  wire n5014_o;
  wire n5015_o;
  wire n5016_o;
  wire n5017_o;
  wire n5018_o;
  wire n5019_o;
  wire n5020_o;
  wire n5021_o;
  wire n5022_o;
  wire n5023_o;
  wire n5024_o;
  wire n5025_o;
  wire n5026_o;
  wire n5027_o;
  wire n5028_o;
  wire n5029_o;
  wire n5030_o;
  wire n5031_o;
  wire n5032_o;
  wire n5033_o;
  wire n5034_o;
  wire n5035_o;
  wire n5036_o;
  wire n5037_o;
  wire n5038_o;
  wire n5039_o;
  wire n5040_o;
  wire n5041_o;
  wire n5042_o;
  wire n5043_o;
  wire n5044_o;
  wire n5045_o;
  wire n5046_o;
  wire n5047_o;
  wire n5048_o;
  wire n5049_o;
  wire n5050_o;
  wire n5051_o;
  wire n5052_o;
  wire n5053_o;
  wire n5054_o;
  wire n5055_o;
  wire n5056_o;
  wire n5057_o;
  wire n5058_o;
  wire n5059_o;
  wire n5060_o;
  wire n5061_o;
  wire n5062_o;
  wire n5063_o;
  wire n5064_o;
  wire n5065_o;
  wire n5066_o;
  wire n5067_o;
  wire n5068_o;
  wire n5069_o;
  wire n5070_o;
  wire n5071_o;
  wire n5072_o;
  wire n5073_o;
  wire n5074_o;
  wire n5075_o;
  wire n5076_o;
  wire n5077_o;
  wire n5078_o;
  wire n5079_o;
  wire n5080_o;
  wire n5081_o;
  wire n5082_o;
  wire n5083_o;
  wire n5084_o;
  wire n5085_o;
  wire n5086_o;
  wire n5087_o;
  wire n5088_o;
  wire n5089_o;
  wire n5090_o;
  wire n5091_o;
  wire n5092_o;
  wire n5093_o;
  wire n5094_o;
  wire n5095_o;
  wire n5096_o;
  wire n5097_o;
  wire n5098_o;
  wire n5099_o;
  wire n5100_o;
  wire n5101_o;
  wire n5102_o;
  wire n5103_o;
  wire n5104_o;
  wire n5105_o;
  wire n5106_o;
  wire n5107_o;
  wire n5108_o;
  wire n5109_o;
  wire n5110_o;
  wire n5111_o;
  wire n5112_o;
  wire n5113_o;
  wire n5114_o;
  wire [10:0] n5117_o;
  wire [41:0] n5118_o;
  wire [41:0] n5123_o;
  wire n5128_o;
  wire n5131_o;
  wire n5132_o;
  wire n5133_o;
  wire n5134_o;
  wire [3:0] n5135_o;
  wire n5137_o;
  wire [3:0] n5138_o;
  wire n5140_o;
  wire n5141_o;
  wire n5142_o;
  wire n5143_o;
  wire n5145_o;
  wire n5146_o;
  wire n5147_o;
  wire n5149_o;
  wire n5150_o;
  wire n5151_o;
  wire [10:0] n5158_o;
  wire n5164_o;
  wire n5166_o;
  wire n5168_o;
  wire n5169_o;
  wire n5170_o;
  wire n5171_o;
  wire n5172_o;
  wire n5173_o;
  wire n5174_o;
  wire n5175_o;
  wire n5176_o;
  wire n5177_o;
  wire n5178_o;
  wire n5179_o;
  wire n5180_o;
  wire n5181_o;
  wire n5182_o;
  wire n5183_o;
  wire n5184_o;
  wire n5185_o;
  wire n5186_o;
  wire n5187_o;
  wire n5188_o;
  wire [18:0] n5192_o;
  wire n5198_o;
  wire n5200_o;
  wire n5202_o;
  wire n5203_o;
  wire n5204_o;
  wire n5205_o;
  wire n5206_o;
  wire n5207_o;
  wire n5208_o;
  wire n5209_o;
  wire n5210_o;
  wire n5211_o;
  wire n5212_o;
  wire n5213_o;
  wire n5214_o;
  wire n5215_o;
  wire n5216_o;
  wire n5217_o;
  wire n5218_o;
  wire n5219_o;
  wire n5220_o;
  wire n5221_o;
  wire n5222_o;
  wire n5223_o;
  wire n5224_o;
  wire n5225_o;
  wire n5226_o;
  wire n5227_o;
  wire n5228_o;
  wire n5229_o;
  wire n5230_o;
  wire n5231_o;
  wire n5232_o;
  wire n5233_o;
  wire n5234_o;
  wire n5235_o;
  wire n5236_o;
  wire n5237_o;
  wire n5238_o;
  wire n5239_o;
  wire n5240_o;
  wire n5241_o;
  wire n5242_o;
  wire n5243_o;
  wire n5244_o;
  wire n5245_o;
  wire n5246_o;
  wire n5247_o;
  wire n5248_o;
  wire n5249_o;
  wire n5250_o;
  wire n5251_o;
  wire n5252_o;
  wire n5253_o;
  wire [30:0] n5255_o;
  wire [31:0] n5257_o;
  wire n5258_o;
  wire [6:0] n5259_o;
  wire n5261_o;
  wire n5262_o;
  wire [31:0] n5263_o;
  wire [30:0] n5264_o;
  wire [31:0] n5266_o;
  wire n5269_o;
  wire n5271_o;
  wire n5273_o;
  wire n5275_o;
  wire n5276_o;
  wire [5:0] n5278_o;
  wire n5279_o;
  wire [6:0] n5280_o;
  wire n5281_o;
  wire n5283_o;
  wire n5285_o;
  wire n5287_o;
  wire n5289_o;
  wire n5291_o;
  wire n5293_o;
  wire n5295_o;
  wire n5297_o;
  wire n5299_o;
  wire n5301_o;
  wire n5303_o;
  wire n5305_o;
  wire n5307_o;
  wire n5309_o;
  wire n5311_o;
  wire n5313_o;
  wire n5315_o;
  wire n5317_o;
  wire n5319_o;
  wire n5321_o;
  wire n5323_o;
  wire n5325_o;
  wire n5327_o;
  wire n5329_o;
  wire n5331_o;
  wire n5333_o;
  wire [6:0] n5337_o;
  wire [6:0] n5338_o;
  wire [6:0] n5339_o;
  wire [6:0] n5340_o;
  wire [6:0] n5341_o;
  wire [6:0] n5342_o;
  wire [6:0] n5343_o;
  wire [6:0] n5344_o;
  wire [6:0] n5345_o;
  wire [6:0] n5346_o;
  wire [6:0] n5347_o;
  wire [6:0] n5348_o;
  wire [6:0] n5349_o;
  wire [6:0] n5350_o;
  wire [6:0] n5351_o;
  wire [6:0] n5352_o;
  wire [6:0] n5353_o;
  wire [6:0] n5354_o;
  wire [6:0] n5355_o;
  wire [6:0] n5356_o;
  wire [6:0] n5357_o;
  wire [6:0] n5358_o;
  wire [6:0] n5359_o;
  wire [6:0] n5360_o;
  wire [6:0] n5361_o;
  wire [6:0] n5362_o;
  wire [6:0] n5363_o;
  wire [6:0] n5364_o;
  wire [6:0] n5365_o;
  wire [6:0] n5366_o;
  wire [6:0] n5367_o;
  wire n5373_o;
  wire [4:0] n5374_o;
  localparam [31:0] n5375_o = 32'b00000000000000000000000000000000;
  wire [26:0] n5376_o;
  wire [31:0] n5377_o;
  wire [31:0] n5378_o;
  wire [1:0] n5379_o;
  wire [31:0] n5380_o;
  wire [31:0] n5381_o;
  wire n5383_o;
  wire [31:0] n5384_o;
  wire [31:0] n5385_o;
  wire [31:0] n5386_o;
  wire n5388_o;
  wire [1:0] n5389_o;
  reg [31:0] n5390_o;
  wire n5393_o;
  wire n5427_o;
  wire n5428_o;
  wire n5429_o;
  wire n5430_o;
  wire n5432_o;
  wire [8:0] n5433_o;
  wire n5435_o;
  wire [2:0] n5436_o;
  wire n5438_o;
  wire n5439_o;
  wire n5440_o;
  wire [1:0] n5441_o;
  wire [1:0] n5442_o;
  wire [1:0] n5443_o;
  wire [2:0] n5444_o;
  wire n5446_o;
  wire n5447_o;
  wire n5448_o;
  wire n5449_o;
  wire [15:0] n5450_o;
  wire [18:0] n5451_o;
  wire [18:0] n5452_o;
  wire [18:0] n5453_o;
  wire [2:0] n5454_o;
  wire n5456_o;
  wire [29:0] n5457_o;
  wire [31:0] n5459_o;
  wire [31:0] n5460_o;
  wire [31:0] n5461_o;
  wire n5466_o;
  wire n5468_o;
  wire n5470_o;
  wire [7:0] n5471_o;
  wire n5473_o;
  wire [3:0] n5474_o;
  wire n5476_o;
  wire [31:0] n5477_o;
  wire [31:0] n5478_o;
  wire [31:0] n5479_o;
  wire [3:0] n5480_o;
  wire n5482_o;
  wire [31:0] n5483_o;
  wire [31:0] n5484_o;
  wire [31:0] n5485_o;
  wire [3:0] n5486_o;
  wire n5488_o;
  wire n5489_o;
  wire [4:0] n5490_o;
  wire [5:0] n5491_o;
  wire [5:0] n5492_o;
  wire [5:0] n5493_o;
  wire [3:0] n5494_o;
  wire n5496_o;
  wire [31:0] n5497_o;
  wire [31:0] n5498_o;
  wire [31:0] n5499_o;
  wire [3:0] n5500_o;
  wire n5502_o;
  wire [15:0] n5503_o;
  wire [15:0] n5504_o;
  wire [37:0] n5505_o;
  wire [63:0] n5506_o;
  wire n5507_o;
  wire [37:0] n5508_o;
  wire [37:0] n5509_o;
  wire [63:0] n5510_o;
  wire [63:0] n5511_o;
  wire [6:0] n5512_o;
  wire n5514_o;
  wire [4:0] n5515_o;
  wire n5517_o;
  wire n5518_o;
  wire n5519_o;
  wire n5520_o;
  wire n5521_o;
  wire n5522_o;
  wire n5523_o;
  wire n5525_o;
  wire n5527_o;
  wire n5528_o;
  wire n5529_o;
  wire [4:0] n5530_o;
  wire [5:0] n5531_o;
  wire [31:0] n5532_o;
  wire [6:0] n5533_o;
  wire [30:0] n5534_o;
  wire [31:0] n5536_o;
  wire n5538_o;
  wire n5540_o;
  wire n5541_o;
  wire n5543_o;
  wire n5545_o;
  wire n5546_o;
  wire n5548_o;
  wire n5549_o;
  wire n5551_o;
  wire n5552_o;
  wire [1:0] n5554_o;
  reg [31:0] n5555_o;
  wire n5558_o;
  wire n5559_o;
  wire n5560_o;
  wire n5563_o;
  wire [2:0] n5565_o;
  wire [2:0] n5566_o;
  wire [2:0] n5567_o;
  wire n5568_o;
  wire n5569_o;
  wire [2:0] n5570_o;
  wire [37:0] n5571_o;
  wire [2:0] n5572_o;
  wire n5573_o;
  wire [37:0] n5574_o;
  wire [37:0] n5575_o;
  wire [31:0] n5576_o;
  wire [31:0] n5577_o;
  wire [34:0] n5578_o;
  wire [133:0] n5579_o;
  wire [1:0] n5580_o;
  wire [1:0] n5581_o;
  wire n5582_o;
  wire n5583_o;
  wire n5584_o;
  wire [18:0] n5585_o;
  wire [34:0] n5586_o;
  wire [34:0] n5587_o;
  wire n5588_o;
  wire n5589_o;
  wire [37:0] n5590_o;
  wire [37:0] n5591_o;
  wire [31:0] n5592_o;
  wire [31:0] n5593_o;
  wire [31:0] n5594_o;
  wire [31:0] n5595_o;
  wire [31:0] n5596_o;
  wire [31:0] n5597_o;
  wire [31:0] n5598_o;
  wire [31:0] n5599_o;
  wire n5601_o;
  wire n5603_o;
  wire [40:0] n5626_o;
  wire [212:0] n5627_o;
  wire [66:0] n5628_o;
  wire [40:0] n5639_o;
  wire [212:0] n5640_o;
  wire [66:0] n5641_o;
  wire n5650_o;
  wire n5651_o;
  localparam [127:0] n5680_o = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam [543:0] n5681_o = 544'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire n5705_o;
  localparam [31:0] n5706_o = 32'b00000000000000000000000000000000;
  wire n5708_o;
  wire n5710_o;
  wire n5712_o;
  wire n5713_o;
  wire n5714_o;
  wire n5715_o;
  wire n5716_o;
  wire [1:0] n5717_o;
  wire n5718_o;
  wire n5719_o;
  wire n5722_o;
  wire n5724_o;
  wire n5741_o;
  wire n5742_o;
  wire n5743_o;
  wire n5744_o;
  wire [15:0] n5745_o;
  wire n5747_o;
  wire [29:0] n5748_o;
  wire [31:0] n5750_o;
  wire n5752_o;
  wire n5754_o;
  wire [31:0] n5755_o;
  wire n5757_o;
  wire [30:0] n5758_o;
  wire [31:0] n5760_o;
  wire n5762_o;
  wire n5763_o;
  wire [4:0] n5764_o;
  wire n5766_o;
  wire [31:0] n5767_o;
  wire n5769_o;
  wire n5770_o;
  wire n5771_o;
  wire n5772_o;
  wire [15:0] n5773_o;
  wire n5775_o;
  wire n5777_o;
  wire n5779_o;
  wire n5780_o;
  wire n5782_o;
  wire n5783_o;
  wire n5785_o;
  wire n5786_o;
  wire n5788_o;
  wire n5790_o;
  wire n5791_o;
  wire n5793_o;
  wire n5794_o;
  wire n5796_o;
  wire n5797_o;
  wire n5799_o;
  wire n5800_o;
  wire n5802_o;
  wire n5803_o;
  wire n5805_o;
  wire n5806_o;
  wire n5808_o;
  wire n5809_o;
  wire n5811_o;
  wire n5812_o;
  wire n5814_o;
  wire n5815_o;
  wire n5817_o;
  wire n5818_o;
  wire n5820_o;
  wire n5821_o;
  wire n5823_o;
  wire n5824_o;
  wire n5826_o;
  wire n5827_o;
  wire n5829_o;
  wire n5830_o;
  wire n5832_o;
  wire n5833_o;
  wire n5834_o;
  wire n5835_o;
  wire n5837_o;
  wire n5839_o;
  wire n5841_o;
  wire n5843_o;
  wire n5845_o;
  wire n5847_o;
  wire n5849_o;
  wire n5851_o;
  wire n5853_o;
  wire n5855_o;
  wire n5857_o;
  wire n5859_o;
  wire n5861_o;
  wire n5863_o;
  wire n5865_o;
  wire n5867_o;
  wire n5869_o;
  wire n5871_o;
  wire n5873_o;
  wire n5875_o;
  wire n5877_o;
  wire n5879_o;
  wire n5881_o;
  wire n5883_o;
  wire n5885_o;
  wire n5887_o;
  wire n5889_o;
  wire n5891_o;
  wire n5893_o;
  wire n5895_o;
  wire [31:0] n5896_o;
  wire n5898_o;
  wire n5900_o;
  wire n5901_o;
  wire [31:0] n5902_o;
  wire n5904_o;
  wire n5906_o;
  wire n5907_o;
  wire [31:0] n5908_o;
  wire n5910_o;
  wire n5912_o;
  wire n5913_o;
  wire n5915_o;
  wire n5917_o;
  wire n5918_o;
  wire n5920_o;
  wire n5922_o;
  wire n5923_o;
  wire n5925_o;
  wire n5927_o;
  wire n5928_o;
  wire n5930_o;
  wire n5932_o;
  wire n5933_o;
  wire n5935_o;
  wire n5937_o;
  wire n5938_o;
  wire n5940_o;
  wire n5942_o;
  wire n5943_o;
  wire n5945_o;
  wire n5947_o;
  wire n5948_o;
  wire n5950_o;
  wire n5952_o;
  wire n5953_o;
  wire n5955_o;
  wire n5957_o;
  wire n5958_o;
  wire n5960_o;
  wire n5962_o;
  wire n5963_o;
  wire n5965_o;
  wire n5967_o;
  wire n5968_o;
  wire n5970_o;
  wire n5972_o;
  wire n5973_o;
  wire n5975_o;
  wire n5977_o;
  wire n5978_o;
  wire n5980_o;
  wire n5982_o;
  wire n5983_o;
  wire n5985_o;
  wire n5987_o;
  wire n5988_o;
  wire n5990_o;
  wire n5992_o;
  wire n5993_o;
  wire n5995_o;
  wire n5997_o;
  wire n5998_o;
  wire n6000_o;
  wire n6002_o;
  wire n6003_o;
  wire n6005_o;
  wire n6007_o;
  wire n6008_o;
  wire n6010_o;
  wire n6012_o;
  wire n6013_o;
  wire n6015_o;
  wire n6017_o;
  wire n6018_o;
  wire n6020_o;
  wire n6022_o;
  wire n6023_o;
  wire n6025_o;
  wire n6027_o;
  wire n6028_o;
  wire n6030_o;
  wire n6032_o;
  wire n6033_o;
  wire n6035_o;
  wire n6037_o;
  wire n6038_o;
  wire n6040_o;
  wire n6042_o;
  wire n6043_o;
  wire n6045_o;
  wire n6047_o;
  wire n6048_o;
  wire n6050_o;
  wire n6052_o;
  wire n6053_o;
  wire n6055_o;
  wire n6057_o;
  wire n6058_o;
  wire [31:0] n6059_o;
  wire n6061_o;
  wire n6063_o;
  wire n6064_o;
  wire [31:0] n6065_o;
  wire n6067_o;
  wire n6069_o;
  wire n6070_o;
  wire [31:0] n6071_o;
  wire n6073_o;
  wire n6075_o;
  wire n6076_o;
  wire n6078_o;
  wire n6080_o;
  wire n6081_o;
  wire n6083_o;
  wire n6085_o;
  wire n6086_o;
  wire n6088_o;
  wire n6090_o;
  wire n6091_o;
  wire n6093_o;
  wire n6095_o;
  wire n6096_o;
  wire n6098_o;
  wire n6100_o;
  wire n6101_o;
  wire n6103_o;
  wire n6105_o;
  wire n6106_o;
  wire n6108_o;
  wire n6110_o;
  wire n6111_o;
  wire n6113_o;
  wire n6115_o;
  wire n6116_o;
  wire n6118_o;
  wire n6120_o;
  wire n6121_o;
  wire n6123_o;
  wire n6125_o;
  wire n6126_o;
  wire n6128_o;
  wire n6130_o;
  wire n6131_o;
  wire n6133_o;
  wire n6135_o;
  wire n6136_o;
  wire n6138_o;
  wire n6140_o;
  wire n6141_o;
  wire n6143_o;
  wire n6145_o;
  wire n6146_o;
  wire n6148_o;
  wire n6150_o;
  wire n6151_o;
  wire n6153_o;
  wire n6155_o;
  wire n6156_o;
  wire n6158_o;
  wire n6160_o;
  wire n6161_o;
  wire n6163_o;
  wire n6165_o;
  wire n6166_o;
  wire n6168_o;
  wire n6170_o;
  wire n6171_o;
  wire n6173_o;
  wire n6175_o;
  wire n6176_o;
  wire n6178_o;
  wire n6180_o;
  wire n6181_o;
  wire n6183_o;
  wire n6185_o;
  wire n6186_o;
  wire n6188_o;
  wire n6190_o;
  wire n6191_o;
  wire n6193_o;
  wire n6195_o;
  wire n6196_o;
  wire n6198_o;
  wire n6200_o;
  wire n6201_o;
  wire n6203_o;
  wire n6205_o;
  wire n6206_o;
  wire n6208_o;
  wire n6210_o;
  wire n6211_o;
  wire n6213_o;
  wire n6215_o;
  wire n6216_o;
  wire n6218_o;
  wire n6220_o;
  wire n6221_o;
  localparam [31:0] n6222_o = 32'b00000000000000000000000000000000;
  wire n6224_o;
  localparam [4:0] n6225_o = 5'b10011;
  wire n6227_o;
  localparam [31:0] n6228_o = 32'b00000001000010000000001100000001;
  wire n6230_o;
  localparam [31:0] n6231_o = 32'b00000000000000000000000000000000;
  wire n6233_o;
  wire n6235_o;
  wire n6237_o;
  wire n6239_o;
  wire n6241_o;
  wire n6243_o;
  wire n6245_o;
  wire n6274_o;
  localparam [31:0] n6275_o = 32'b00000000000000000000000000000000;
  wire [119:0] n6276_o;
  wire n6277_o;
  wire n6278_o;
  wire n6279_o;
  wire n6280_o;
  wire n6281_o;
  wire n6282_o;
  wire n6283_o;
  wire n6284_o;
  wire n6285_o;
  wire n6286_o;
  wire n6287_o;
  wire n6288_o;
  wire n6289_o;
  wire n6290_o;
  wire n6291_o;
  wire n6292_o;
  wire n6293_o;
  reg n6294_o;
  wire n6295_o;
  wire n6296_o;
  wire n6297_o;
  wire n6298_o;
  wire n6299_o;
  wire n6300_o;
  wire n6301_o;
  wire n6302_o;
  wire n6303_o;
  wire n6304_o;
  wire n6305_o;
  wire n6306_o;
  wire n6307_o;
  wire n6308_o;
  wire n6309_o;
  wire n6310_o;
  wire n6311_o;
  reg n6312_o;
  wire n6313_o;
  wire n6314_o;
  wire n6315_o;
  wire n6316_o;
  wire n6317_o;
  wire n6318_o;
  wire n6319_o;
  wire n6320_o;
  wire n6321_o;
  wire n6322_o;
  wire n6323_o;
  wire n6324_o;
  wire n6325_o;
  wire n6326_o;
  wire n6327_o;
  wire n6328_o;
  wire n6329_o;
  reg n6330_o;
  wire n6331_o;
  wire n6332_o;
  wire n6333_o;
  wire n6334_o;
  wire n6335_o;
  wire n6336_o;
  wire n6337_o;
  wire n6338_o;
  wire n6339_o;
  wire n6340_o;
  wire n6341_o;
  wire n6342_o;
  wire n6343_o;
  wire n6344_o;
  wire n6345_o;
  wire n6346_o;
  wire n6347_o;
  reg n6348_o;
  wire n6349_o;
  wire n6350_o;
  wire n6351_o;
  wire n6352_o;
  wire n6353_o;
  wire n6354_o;
  wire n6355_o;
  wire n6356_o;
  wire n6357_o;
  wire n6358_o;
  wire n6359_o;
  wire n6360_o;
  wire n6361_o;
  wire n6362_o;
  wire n6363_o;
  wire n6364_o;
  wire n6365_o;
  reg n6366_o;
  wire n6367_o;
  wire n6368_o;
  wire n6369_o;
  wire n6370_o;
  wire n6371_o;
  wire n6372_o;
  wire n6373_o;
  wire n6374_o;
  wire n6375_o;
  wire n6376_o;
  wire n6377_o;
  wire n6378_o;
  wire n6379_o;
  wire n6380_o;
  wire n6381_o;
  reg n6382_o;
  wire n6383_o;
  wire n6384_o;
  wire n6385_o;
  wire n6386_o;
  wire n6387_o;
  wire n6388_o;
  wire n6389_o;
  wire n6390_o;
  wire n6391_o;
  wire n6392_o;
  wire n6393_o;
  wire n6394_o;
  wire n6395_o;
  wire n6396_o;
  wire n6397_o;
  reg n6398_o;
  wire n6399_o;
  wire n6400_o;
  wire n6401_o;
  wire n6402_o;
  wire n6403_o;
  wire n6404_o;
  wire n6405_o;
  wire n6406_o;
  wire n6407_o;
  wire n6408_o;
  wire n6409_o;
  wire n6410_o;
  wire n6411_o;
  wire n6412_o;
  wire n6413_o;
  reg n6414_o;
  wire n6415_o;
  wire n6416_o;
  wire n6417_o;
  wire n6418_o;
  wire n6419_o;
  wire n6420_o;
  wire n6421_o;
  wire n6422_o;
  wire n6423_o;
  wire n6424_o;
  wire n6425_o;
  wire n6426_o;
  wire n6427_o;
  wire n6428_o;
  wire n6429_o;
  reg n6430_o;
  wire n6431_o;
  wire n6432_o;
  wire n6433_o;
  wire n6434_o;
  wire n6435_o;
  wire n6436_o;
  wire n6437_o;
  wire n6438_o;
  wire n6439_o;
  wire n6440_o;
  wire n6441_o;
  wire n6442_o;
  wire n6443_o;
  wire n6444_o;
  wire n6445_o;
  reg n6446_o;
  wire n6447_o;
  wire n6448_o;
  wire n6449_o;
  wire n6450_o;
  wire n6451_o;
  wire n6452_o;
  wire n6453_o;
  wire n6454_o;
  wire n6455_o;
  wire n6456_o;
  wire n6457_o;
  wire n6458_o;
  wire n6459_o;
  wire n6460_o;
  wire n6461_o;
  reg n6462_o;
  wire n6463_o;
  wire n6464_o;
  wire n6465_o;
  wire n6466_o;
  wire n6467_o;
  wire n6468_o;
  wire n6469_o;
  wire n6470_o;
  wire n6471_o;
  wire n6472_o;
  wire n6473_o;
  wire n6474_o;
  wire n6475_o;
  wire n6476_o;
  wire n6477_o;
  wire n6478_o;
  reg n6479_o;
  wire n6480_o;
  wire n6481_o;
  wire n6482_o;
  wire n6483_o;
  wire n6484_o;
  wire n6485_o;
  wire n6486_o;
  wire n6487_o;
  wire n6488_o;
  wire n6489_o;
  wire n6490_o;
  wire n6491_o;
  wire n6492_o;
  wire n6493_o;
  wire n6494_o;
  wire n6495_o;
  reg n6496_o;
  wire [2:0] n6497_o;
  wire [2:0] n6498_o;
  wire [2:0] n6499_o;
  wire [2:0] n6500_o;
  wire [2:0] n6501_o;
  wire [2:0] n6502_o;
  wire [2:0] n6503_o;
  wire [2:0] n6504_o;
  wire [2:0] n6505_o;
  wire [2:0] n6506_o;
  wire [2:0] n6507_o;
  wire [2:0] n6508_o;
  wire [2:0] n6509_o;
  wire [2:0] n6510_o;
  wire [2:0] n6511_o;
  reg [2:0] n6512_o;
  wire n6513_o;
  wire n6514_o;
  wire n6515_o;
  wire n6516_o;
  wire n6517_o;
  wire n6518_o;
  wire n6519_o;
  wire n6520_o;
  wire n6521_o;
  wire n6522_o;
  wire n6523_o;
  wire n6524_o;
  wire n6525_o;
  wire n6526_o;
  wire n6527_o;
  wire n6528_o;
  wire n6529_o;
  reg n6530_o;
  wire n6531_o;
  wire n6532_o;
  wire n6533_o;
  wire n6534_o;
  wire n6535_o;
  wire n6536_o;
  wire n6537_o;
  wire n6538_o;
  wire n6539_o;
  wire n6540_o;
  wire n6541_o;
  wire n6542_o;
  wire n6543_o;
  wire n6544_o;
  wire n6545_o;
  wire n6546_o;
  wire n6547_o;
  reg n6548_o;
  wire [1:0] n6549_o;
  wire [1:0] n6550_o;
  wire [1:0] n6551_o;
  wire [1:0] n6552_o;
  wire [1:0] n6553_o;
  wire [1:0] n6554_o;
  wire [1:0] n6555_o;
  wire [1:0] n6556_o;
  wire [1:0] n6557_o;
  wire [1:0] n6558_o;
  wire [1:0] n6559_o;
  wire [1:0] n6560_o;
  wire [1:0] n6561_o;
  wire [1:0] n6562_o;
  wire [1:0] n6563_o;
  wire [1:0] n6564_o;
  wire [1:0] n6565_o;
  reg [1:0] n6566_o;
  wire n6567_o;
  wire n6568_o;
  wire n6569_o;
  wire n6570_o;
  wire n6571_o;
  wire n6572_o;
  wire n6573_o;
  wire n6574_o;
  wire n6575_o;
  wire n6576_o;
  wire n6577_o;
  wire n6578_o;
  wire n6579_o;
  wire n6580_o;
  wire n6581_o;
  wire n6582_o;
  wire n6583_o;
  reg n6584_o;
  wire n6585_o;
  wire n6586_o;
  wire n6587_o;
  wire n6588_o;
  wire n6589_o;
  wire n6590_o;
  wire n6591_o;
  wire n6592_o;
  wire n6593_o;
  wire n6594_o;
  wire n6595_o;
  wire n6596_o;
  wire n6597_o;
  wire n6598_o;
  wire n6599_o;
  wire n6600_o;
  wire n6601_o;
  reg n6602_o;
  wire n6603_o;
  wire n6604_o;
  wire n6605_o;
  wire n6606_o;
  wire n6607_o;
  wire n6608_o;
  wire n6609_o;
  wire n6610_o;
  wire n6611_o;
  wire n6612_o;
  wire n6613_o;
  wire n6614_o;
  wire n6615_o;
  wire n6616_o;
  wire n6617_o;
  wire n6618_o;
  wire n6619_o;
  reg n6620_o;
  wire n6621_o;
  wire n6622_o;
  wire n6623_o;
  wire n6624_o;
  wire n6625_o;
  wire n6626_o;
  wire n6627_o;
  wire n6628_o;
  wire n6629_o;
  wire n6630_o;
  wire n6631_o;
  wire n6632_o;
  wire n6633_o;
  wire n6634_o;
  wire n6635_o;
  wire n6636_o;
  wire n6637_o;
  reg n6638_o;
  wire [5:0] n6639_o;
  wire [5:0] n6640_o;
  wire [5:0] n6641_o;
  wire [5:0] n6642_o;
  wire [5:0] n6643_o;
  wire [5:0] n6644_o;
  wire [5:0] n6645_o;
  wire [5:0] n6646_o;
  wire [5:0] n6647_o;
  wire [5:0] n6648_o;
  wire [5:0] n6649_o;
  wire [5:0] n6650_o;
  wire [5:0] n6651_o;
  wire [5:0] n6652_o;
  wire [5:0] n6653_o;
  wire [5:0] n6654_o;
  wire [5:0] n6655_o;
  reg [5:0] n6656_o;
  wire n6657_o;
  wire n6658_o;
  wire n6659_o;
  wire n6660_o;
  wire n6661_o;
  wire n6662_o;
  wire n6663_o;
  wire n6664_o;
  wire n6665_o;
  wire n6666_o;
  wire n6667_o;
  wire n6668_o;
  wire n6669_o;
  wire n6670_o;
  wire n6671_o;
  wire n6672_o;
  wire n6673_o;
  reg n6674_o;
  wire n6675_o;
  wire n6676_o;
  wire n6677_o;
  wire n6678_o;
  wire n6679_o;
  wire n6680_o;
  wire n6681_o;
  wire n6682_o;
  wire n6683_o;
  wire n6684_o;
  wire n6685_o;
  wire n6686_o;
  wire n6687_o;
  wire n6688_o;
  wire n6689_o;
  wire n6690_o;
  wire n6691_o;
  reg n6692_o;
  wire [31:0] n6716_o;
  wire [1:0] n6722_o;
  wire n6723_o;
  wire [2:0] n6724_o;
  wire n6725_o;
  wire [3:0] n6726_o;
  wire [7:0] n6727_o;
  wire [11:0] n6728_o;
  wire n6729_o;
  wire [11:0] n6730_o;
  wire [31:0] n6732_o;
  localparam [31:0] n6734_o = 32'b00000000000000000000000000000000;
  localparam [31:0] n6735_o = 32'b00000000000000000000000000000000;
  wire n6736_o;
  wire [3:0] n6737_o;
  wire n6739_o;
  wire n6740_o;
  wire n6741_o;
  wire n6742_o;
  wire [4:0] n6743_o;
  wire [4:0] n6748_o;
  wire [31:0] n6753_o;
  wire [31:0] n6754_o;
  wire [63:0] n6755_o;
  wire [63:0] n6756_o;
  wire [63:0] n6757_o;
  wire n6760_o;
  wire n6765_o;
  wire [31:0] n6766_o;
  wire [31:0] n6767_o;
  wire [31:0] n6768_o;
  wire n6769_o;
  wire n6770_o;
  wire [31:0] n6771_o;
  wire [31:0] n6772_o;
  wire n6773_o;
  wire [31:0] n6774_o;
  wire [31:0] n6775_o;
  wire [31:0] n6776_o;
  wire [31:0] n6787_o;
  wire [32:0] n6789_o;
  wire [32:0] n6791_o;
  wire n6792_o;
  wire [32:0] n6793_o;
  wire [31:0] n6794_o;
  wire [32:0] n6796_o;
  wire [32:0] n6798_o;
  wire n6800_o;
  wire n6805_o;
  wire [31:0] n6806_o;
  wire [31:0] n6807_o;
  wire [31:0] n6808_o;
  wire n6809_o;
  wire n6810_o;
  wire [31:0] n6811_o;
  wire [31:0] n6812_o;
  wire n6813_o;
  wire [31:0] n6814_o;
  wire [31:0] n6815_o;
  wire [31:0] n6816_o;
  wire [31:0] n6827_o;
  wire [32:0] n6829_o;
  wire [32:0] n6831_o;
  wire n6832_o;
  wire [32:0] n6833_o;
  wire [31:0] n6834_o;
  wire [32:0] n6836_o;
  wire [32:0] n6838_o;
  wire n6840_o;
  wire n6845_o;
  wire [31:0] n6846_o;
  wire [31:0] n6847_o;
  wire [31:0] n6848_o;
  wire n6849_o;
  wire n6850_o;
  wire [31:0] n6851_o;
  wire [31:0] n6852_o;
  wire n6853_o;
  wire [31:0] n6854_o;
  wire [31:0] n6855_o;
  wire [31:0] n6856_o;
  wire [31:0] n6867_o;
  wire [32:0] n6869_o;
  wire [32:0] n6871_o;
  wire n6872_o;
  wire [32:0] n6873_o;
  wire [31:0] n6874_o;
  wire [32:0] n6876_o;
  wire [32:0] n6878_o;
  wire n6880_o;
  wire n6885_o;
  wire [31:0] n6886_o;
  wire [31:0] n6887_o;
  wire [31:0] n6888_o;
  wire n6889_o;
  wire n6890_o;
  wire [31:0] n6891_o;
  wire [31:0] n6892_o;
  wire n6893_o;
  wire [31:0] n6894_o;
  wire [31:0] n6895_o;
  wire [31:0] n6896_o;
  wire [31:0] n6907_o;
  wire [32:0] n6909_o;
  wire [32:0] n6911_o;
  wire n6912_o;
  wire [32:0] n6913_o;
  wire [31:0] n6914_o;
  wire [32:0] n6916_o;
  wire [32:0] n6918_o;
  wire n6920_o;
  wire n6925_o;
  wire [31:0] n6926_o;
  wire [31:0] n6927_o;
  wire [31:0] n6928_o;
  wire n6929_o;
  wire n6930_o;
  wire [31:0] n6931_o;
  wire [31:0] n6932_o;
  wire n6933_o;
  wire [31:0] n6934_o;
  wire [31:0] n6935_o;
  wire [31:0] n6936_o;
  wire [31:0] n6947_o;
  wire [32:0] n6949_o;
  wire [32:0] n6951_o;
  wire n6952_o;
  wire [32:0] n6953_o;
  wire [31:0] n6954_o;
  wire [32:0] n6956_o;
  wire [32:0] n6958_o;
  wire n6960_o;
  wire n6965_o;
  wire [31:0] n6966_o;
  wire [31:0] n6967_o;
  wire [31:0] n6968_o;
  wire n6969_o;
  wire n6970_o;
  wire [31:0] n6971_o;
  wire [31:0] n6972_o;
  wire n6973_o;
  wire [31:0] n6974_o;
  wire [31:0] n6975_o;
  wire [31:0] n6976_o;
  wire [31:0] n6987_o;
  wire [32:0] n6989_o;
  wire [32:0] n6991_o;
  wire n6992_o;
  wire [32:0] n6993_o;
  wire [31:0] n6994_o;
  wire [32:0] n6996_o;
  wire [32:0] n6998_o;
  wire n7000_o;
  wire n7005_o;
  wire [31:0] n7006_o;
  wire [31:0] n7007_o;
  wire [31:0] n7008_o;
  wire n7009_o;
  wire n7010_o;
  wire [31:0] n7011_o;
  wire [31:0] n7012_o;
  wire n7013_o;
  wire [31:0] n7014_o;
  wire [31:0] n7015_o;
  wire [31:0] n7016_o;
  wire [31:0] n7027_o;
  wire [32:0] n7029_o;
  wire [32:0] n7031_o;
  wire n7032_o;
  wire [32:0] n7033_o;
  wire [31:0] n7034_o;
  wire [32:0] n7036_o;
  wire [32:0] n7038_o;
  wire n7040_o;
  wire n7045_o;
  wire [31:0] n7046_o;
  wire [31:0] n7047_o;
  wire [31:0] n7048_o;
  wire n7049_o;
  wire n7050_o;
  wire [31:0] n7051_o;
  wire [31:0] n7052_o;
  wire n7053_o;
  wire [31:0] n7054_o;
  wire [31:0] n7055_o;
  wire [31:0] n7056_o;
  wire [31:0] n7067_o;
  wire [32:0] n7069_o;
  wire [32:0] n7071_o;
  wire n7072_o;
  wire [32:0] n7073_o;
  wire [31:0] n7074_o;
  wire [32:0] n7076_o;
  wire [32:0] n7078_o;
  wire n7080_o;
  wire n7085_o;
  wire [31:0] n7086_o;
  wire [31:0] n7087_o;
  wire [31:0] n7088_o;
  wire n7089_o;
  wire n7090_o;
  wire [31:0] n7091_o;
  wire [31:0] n7092_o;
  wire n7093_o;
  wire [31:0] n7094_o;
  wire [31:0] n7095_o;
  wire [31:0] n7096_o;
  wire [31:0] n7107_o;
  wire [32:0] n7109_o;
  wire [32:0] n7111_o;
  wire n7112_o;
  wire [32:0] n7113_o;
  wire [31:0] n7114_o;
  wire [32:0] n7116_o;
  wire [32:0] n7118_o;
  wire n7120_o;
  wire n7125_o;
  wire [31:0] n7126_o;
  wire [31:0] n7127_o;
  wire [31:0] n7128_o;
  wire n7129_o;
  wire n7130_o;
  wire [31:0] n7131_o;
  wire [31:0] n7132_o;
  wire n7133_o;
  wire [31:0] n7134_o;
  wire [31:0] n7135_o;
  wire [31:0] n7136_o;
  wire [31:0] n7147_o;
  wire [32:0] n7149_o;
  wire [32:0] n7151_o;
  wire n7152_o;
  wire [32:0] n7153_o;
  wire [31:0] n7154_o;
  wire [32:0] n7156_o;
  wire [32:0] n7158_o;
  wire n7160_o;
  wire n7165_o;
  wire [31:0] n7166_o;
  wire [31:0] n7167_o;
  wire [31:0] n7168_o;
  wire n7169_o;
  wire n7170_o;
  wire [31:0] n7171_o;
  wire [31:0] n7172_o;
  wire n7173_o;
  wire [31:0] n7174_o;
  wire [31:0] n7175_o;
  wire [31:0] n7176_o;
  wire [31:0] n7187_o;
  wire [32:0] n7189_o;
  wire [32:0] n7191_o;
  wire n7192_o;
  wire [32:0] n7193_o;
  wire [31:0] n7194_o;
  wire [32:0] n7196_o;
  wire [32:0] n7198_o;
  wire n7200_o;
  wire n7205_o;
  wire [31:0] n7206_o;
  wire [31:0] n7207_o;
  wire [31:0] n7208_o;
  wire n7209_o;
  wire n7210_o;
  wire [31:0] n7211_o;
  wire [31:0] n7212_o;
  wire n7213_o;
  wire [31:0] n7214_o;
  wire [31:0] n7215_o;
  wire [31:0] n7216_o;
  wire [31:0] n7227_o;
  wire [32:0] n7229_o;
  wire [32:0] n7231_o;
  wire n7232_o;
  wire [32:0] n7233_o;
  wire [31:0] n7234_o;
  wire [32:0] n7236_o;
  wire [32:0] n7238_o;
  wire n7240_o;
  wire n7245_o;
  wire [31:0] n7246_o;
  wire [31:0] n7247_o;
  wire [31:0] n7248_o;
  wire n7249_o;
  wire n7250_o;
  wire [31:0] n7251_o;
  wire [31:0] n7252_o;
  wire n7253_o;
  wire [31:0] n7254_o;
  wire [31:0] n7255_o;
  wire [31:0] n7256_o;
  wire [31:0] n7267_o;
  wire [32:0] n7269_o;
  wire [32:0] n7271_o;
  wire n7272_o;
  wire [32:0] n7273_o;
  wire [31:0] n7274_o;
  wire [32:0] n7276_o;
  wire [32:0] n7278_o;
  wire n7280_o;
  wire n7285_o;
  wire [31:0] n7286_o;
  wire [31:0] n7287_o;
  wire [31:0] n7288_o;
  wire n7289_o;
  wire n7290_o;
  wire [31:0] n7291_o;
  wire [31:0] n7292_o;
  wire n7293_o;
  wire [31:0] n7294_o;
  wire [31:0] n7295_o;
  wire [31:0] n7296_o;
  wire [31:0] n7307_o;
  wire [32:0] n7309_o;
  wire [32:0] n7311_o;
  wire n7312_o;
  wire [32:0] n7313_o;
  wire [31:0] n7314_o;
  wire [32:0] n7316_o;
  wire [32:0] n7318_o;
  wire n7320_o;
  wire n7325_o;
  wire [31:0] n7326_o;
  wire [31:0] n7327_o;
  wire [31:0] n7328_o;
  wire n7329_o;
  wire n7330_o;
  wire [31:0] n7331_o;
  wire [31:0] n7332_o;
  wire n7333_o;
  wire [31:0] n7334_o;
  wire [31:0] n7335_o;
  wire [31:0] n7336_o;
  wire [31:0] n7347_o;
  wire [32:0] n7349_o;
  wire [32:0] n7351_o;
  wire n7352_o;
  wire [32:0] n7353_o;
  wire [31:0] n7354_o;
  wire [32:0] n7356_o;
  wire [32:0] n7358_o;
  wire n7360_o;
  wire n7365_o;
  wire [31:0] n7366_o;
  wire [31:0] n7367_o;
  wire [31:0] n7368_o;
  wire n7369_o;
  wire n7370_o;
  wire [31:0] n7371_o;
  wire [31:0] n7372_o;
  wire n7373_o;
  wire [31:0] n7374_o;
  wire [31:0] n7375_o;
  wire [31:0] n7376_o;
  wire [31:0] n7387_o;
  wire [32:0] n7389_o;
  wire [32:0] n7391_o;
  wire n7392_o;
  wire [32:0] n7393_o;
  wire [31:0] n7394_o;
  wire [32:0] n7396_o;
  wire [32:0] n7398_o;
  wire n7400_o;
  wire n7405_o;
  wire [31:0] n7406_o;
  wire [31:0] n7407_o;
  wire [31:0] n7408_o;
  wire n7409_o;
  wire n7410_o;
  wire [31:0] n7411_o;
  wire [31:0] n7412_o;
  wire n7413_o;
  wire [31:0] n7414_o;
  wire [31:0] n7415_o;
  wire [31:0] n7416_o;
  wire [31:0] n7427_o;
  wire [32:0] n7429_o;
  wire [32:0] n7431_o;
  wire n7432_o;
  wire [32:0] n7433_o;
  wire [31:0] n7434_o;
  wire [32:0] n7436_o;
  wire [32:0] n7438_o;
  wire n7440_o;
  wire n7445_o;
  wire [31:0] n7446_o;
  wire [31:0] n7447_o;
  wire [31:0] n7448_o;
  wire n7449_o;
  wire n7450_o;
  wire [31:0] n7451_o;
  wire [31:0] n7452_o;
  wire n7453_o;
  wire [31:0] n7454_o;
  wire [31:0] n7455_o;
  wire [31:0] n7456_o;
  wire [31:0] n7467_o;
  wire [32:0] n7469_o;
  wire [32:0] n7471_o;
  wire n7472_o;
  wire [32:0] n7473_o;
  wire [31:0] n7474_o;
  wire [32:0] n7476_o;
  wire [32:0] n7478_o;
  wire n7480_o;
  wire n7485_o;
  wire [31:0] n7486_o;
  wire [31:0] n7487_o;
  wire [31:0] n7488_o;
  wire n7489_o;
  wire n7490_o;
  wire [31:0] n7491_o;
  wire [31:0] n7492_o;
  wire n7493_o;
  wire [31:0] n7494_o;
  wire [31:0] n7495_o;
  wire [31:0] n7496_o;
  wire [31:0] n7507_o;
  wire [32:0] n7509_o;
  wire [32:0] n7511_o;
  wire n7512_o;
  wire [32:0] n7513_o;
  wire [31:0] n7514_o;
  wire [32:0] n7516_o;
  wire [32:0] n7518_o;
  wire n7520_o;
  wire n7525_o;
  wire [31:0] n7526_o;
  wire [31:0] n7527_o;
  wire [31:0] n7528_o;
  wire n7529_o;
  wire n7530_o;
  wire [31:0] n7531_o;
  wire [31:0] n7532_o;
  wire n7533_o;
  wire [31:0] n7534_o;
  wire [31:0] n7535_o;
  wire [31:0] n7536_o;
  wire [31:0] n7547_o;
  wire [32:0] n7549_o;
  wire [32:0] n7551_o;
  wire n7552_o;
  wire [32:0] n7553_o;
  wire [31:0] n7554_o;
  wire [32:0] n7556_o;
  wire [32:0] n7558_o;
  wire n7560_o;
  wire n7565_o;
  wire [31:0] n7566_o;
  wire [31:0] n7567_o;
  wire [31:0] n7568_o;
  wire n7569_o;
  wire n7570_o;
  wire [31:0] n7571_o;
  wire [31:0] n7572_o;
  wire n7573_o;
  wire [31:0] n7574_o;
  wire [31:0] n7575_o;
  wire [31:0] n7576_o;
  wire [31:0] n7587_o;
  wire [32:0] n7589_o;
  wire [32:0] n7591_o;
  wire n7592_o;
  wire [32:0] n7593_o;
  wire [31:0] n7594_o;
  wire [32:0] n7596_o;
  wire [32:0] n7598_o;
  wire n7600_o;
  wire n7605_o;
  wire [31:0] n7606_o;
  wire [31:0] n7607_o;
  wire [31:0] n7608_o;
  wire n7609_o;
  wire n7610_o;
  wire [31:0] n7611_o;
  wire [31:0] n7612_o;
  wire n7613_o;
  wire [31:0] n7614_o;
  wire [31:0] n7615_o;
  wire [31:0] n7616_o;
  wire [31:0] n7627_o;
  wire [32:0] n7629_o;
  wire [32:0] n7631_o;
  wire n7632_o;
  wire [32:0] n7633_o;
  wire [31:0] n7634_o;
  wire [32:0] n7636_o;
  wire [32:0] n7638_o;
  wire n7640_o;
  wire n7645_o;
  wire [31:0] n7646_o;
  wire [31:0] n7647_o;
  wire [31:0] n7648_o;
  wire n7649_o;
  wire n7650_o;
  wire [31:0] n7651_o;
  wire [31:0] n7652_o;
  wire n7653_o;
  wire [31:0] n7654_o;
  wire [31:0] n7655_o;
  wire [31:0] n7656_o;
  wire [31:0] n7667_o;
  wire [32:0] n7669_o;
  wire [32:0] n7671_o;
  wire n7672_o;
  wire [32:0] n7673_o;
  wire [31:0] n7674_o;
  wire [32:0] n7676_o;
  wire [32:0] n7678_o;
  wire n7680_o;
  wire n7685_o;
  wire [31:0] n7686_o;
  wire [31:0] n7687_o;
  wire [31:0] n7688_o;
  wire n7689_o;
  wire n7690_o;
  wire [31:0] n7691_o;
  wire [31:0] n7692_o;
  wire n7693_o;
  wire [31:0] n7694_o;
  wire [31:0] n7695_o;
  wire [31:0] n7696_o;
  wire [31:0] n7707_o;
  wire [32:0] n7709_o;
  wire [32:0] n7711_o;
  wire n7712_o;
  wire [32:0] n7713_o;
  wire [31:0] n7714_o;
  wire [32:0] n7716_o;
  wire [32:0] n7718_o;
  wire n7720_o;
  wire n7725_o;
  wire [31:0] n7726_o;
  wire [31:0] n7727_o;
  wire [31:0] n7728_o;
  wire n7729_o;
  wire n7730_o;
  wire [31:0] n7731_o;
  wire [31:0] n7732_o;
  wire n7733_o;
  wire [31:0] n7734_o;
  wire [31:0] n7735_o;
  wire [31:0] n7736_o;
  wire [31:0] n7747_o;
  wire [32:0] n7749_o;
  wire [32:0] n7751_o;
  wire n7752_o;
  wire [32:0] n7753_o;
  wire [31:0] n7754_o;
  wire [32:0] n7756_o;
  wire [32:0] n7758_o;
  wire n7760_o;
  wire n7765_o;
  wire [31:0] n7766_o;
  wire [31:0] n7767_o;
  wire [31:0] n7768_o;
  wire n7769_o;
  wire n7770_o;
  wire [31:0] n7771_o;
  wire [31:0] n7772_o;
  wire n7773_o;
  wire [31:0] n7774_o;
  wire [31:0] n7775_o;
  wire [31:0] n7776_o;
  wire [31:0] n7787_o;
  wire [32:0] n7789_o;
  wire [32:0] n7791_o;
  wire n7792_o;
  wire [32:0] n7793_o;
  wire [31:0] n7794_o;
  wire [32:0] n7796_o;
  wire [32:0] n7798_o;
  wire n7800_o;
  wire n7805_o;
  wire [31:0] n7806_o;
  wire [31:0] n7807_o;
  wire [31:0] n7808_o;
  wire n7809_o;
  wire n7810_o;
  wire [31:0] n7811_o;
  wire [31:0] n7812_o;
  wire n7813_o;
  wire [31:0] n7814_o;
  wire [31:0] n7815_o;
  wire [31:0] n7816_o;
  wire [31:0] n7827_o;
  wire [32:0] n7829_o;
  wire [32:0] n7831_o;
  wire n7832_o;
  wire [32:0] n7833_o;
  wire [31:0] n7834_o;
  wire [32:0] n7836_o;
  wire [32:0] n7838_o;
  wire n7840_o;
  wire n7845_o;
  wire [31:0] n7846_o;
  wire [31:0] n7847_o;
  wire [31:0] n7848_o;
  wire n7849_o;
  wire n7850_o;
  wire [31:0] n7851_o;
  wire [31:0] n7852_o;
  wire n7853_o;
  wire [31:0] n7854_o;
  wire [31:0] n7855_o;
  wire [31:0] n7856_o;
  wire [31:0] n7867_o;
  wire [32:0] n7869_o;
  wire [32:0] n7871_o;
  wire n7872_o;
  wire [32:0] n7873_o;
  wire [31:0] n7874_o;
  wire [32:0] n7876_o;
  wire [32:0] n7878_o;
  wire n7880_o;
  wire n7885_o;
  wire [31:0] n7886_o;
  wire [31:0] n7887_o;
  wire [31:0] n7888_o;
  wire n7889_o;
  wire n7890_o;
  wire [31:0] n7891_o;
  wire [31:0] n7892_o;
  wire n7893_o;
  wire [31:0] n7894_o;
  wire [31:0] n7895_o;
  wire [31:0] n7896_o;
  wire [31:0] n7907_o;
  wire [32:0] n7909_o;
  wire [32:0] n7911_o;
  wire n7912_o;
  wire [32:0] n7913_o;
  wire [31:0] n7914_o;
  wire [32:0] n7916_o;
  wire [32:0] n7918_o;
  wire n7920_o;
  wire n7925_o;
  wire [31:0] n7926_o;
  wire [31:0] n7927_o;
  wire [31:0] n7928_o;
  wire n7929_o;
  wire n7930_o;
  wire [31:0] n7931_o;
  wire [31:0] n7932_o;
  wire n7933_o;
  wire [31:0] n7934_o;
  wire [31:0] n7935_o;
  wire [31:0] n7936_o;
  wire [31:0] n7947_o;
  wire [32:0] n7949_o;
  wire [32:0] n7951_o;
  wire n7952_o;
  wire [32:0] n7953_o;
  wire [31:0] n7954_o;
  wire [32:0] n7956_o;
  wire [32:0] n7958_o;
  wire n7960_o;
  wire n7965_o;
  wire [31:0] n7966_o;
  wire [31:0] n7967_o;
  wire [31:0] n7968_o;
  wire n7969_o;
  wire n7970_o;
  wire [31:0] n7971_o;
  wire [31:0] n7972_o;
  wire n7973_o;
  wire [31:0] n7974_o;
  wire [31:0] n7975_o;
  wire [31:0] n7976_o;
  wire [31:0] n7987_o;
  wire [32:0] n7989_o;
  wire [32:0] n7991_o;
  wire n7992_o;
  wire [32:0] n7993_o;
  wire [31:0] n7994_o;
  wire [32:0] n7996_o;
  wire [32:0] n7998_o;
  wire n8000_o;
  wire n8005_o;
  wire [31:0] n8006_o;
  wire [31:0] n8007_o;
  wire [31:0] n8008_o;
  wire n8009_o;
  wire n8010_o;
  wire [31:0] n8011_o;
  wire [31:0] n8012_o;
  wire n8013_o;
  wire [31:0] n8014_o;
  wire [31:0] n8015_o;
  wire [31:0] n8016_o;
  wire [31:0] n8027_o;
  wire [32:0] n8029_o;
  wire [32:0] n8031_o;
  wire n8032_o;
  wire [32:0] n8033_o;
  wire [31:0] n8034_o;
  wire [32:0] n8036_o;
  wire [32:0] n8038_o;
  wire [31:0] n8040_o;
  localparam [1023:0] n8041_o = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire [31:0] n8043_o;
  localparam [1023:0] n8044_o = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire [31:0] n8046_o;
  wire [31:0] n8048_o;
  wire [31:0] n8050_o;
  wire [927:0] n8051_o;
  wire [31:0] n8052_o;
  wire [927:0] n8053_o;
  localparam [31:0] n8057_o = 32'b00000000000000000000000000000000;
  wire n8058_o;
  wire n8059_o;
  wire n8060_o;
  wire n8061_o;
  wire n8062_o;
  wire n8063_o;
  wire n8064_o;
  wire n8066_o;
  wire n8067_o;
  wire n8068_o;
  wire n8069_o;
  wire n8070_o;
  wire n8071_o;
  wire n8072_o;
  wire n8074_o;
  wire n8075_o;
  wire n8076_o;
  wire n8077_o;
  wire n8078_o;
  wire n8079_o;
  wire n8080_o;
  wire [28:0] n8081_o;
  wire [31:0] n8082_o;
  wire n8087_o;
  wire n8088_o;
  wire n8089_o;
  wire [3:0] n8093_o;
  wire n8095_o;
  wire n8096_o;
  wire [3:0] n8099_o;
  wire n8101_o;
  wire n8102_o;
  wire n8103_o;
  wire n8104_o;
  wire [1:0] n8107_o;
  wire n8109_o;
  wire [1:0] n8110_o;
  wire n8112_o;
  wire n8113_o;
  wire n8114_o;
  wire [3:0] n8117_o;
  wire n8119_o;
  wire [3:0] n8120_o;
  wire n8122_o;
  wire n8123_o;
  wire n8124_o;
  wire [3:0] n8127_o;
  wire n8129_o;
  wire n8130_o;
  wire n8133_o;
  wire n8134_o;
  wire n8135_o;
  wire n8136_o;
  wire n8137_o;
  wire n8140_o;
  wire n8141_o;
  wire n8142_o;
  wire n8143_o;
  wire [3:0] n8146_o;
  wire n8148_o;
  wire [3:0] n8149_o;
  wire n8151_o;
  wire n8152_o;
  wire n8153_o;
  wire [3:0] n8156_o;
  wire n8158_o;
  wire n8159_o;
  wire n8160_o;
  wire n8161_o;
  wire [3:0] n8164_o;
  wire n8166_o;
  wire n8167_o;
  wire n8168_o;
  wire n8169_o;
  wire n8170_o;
  wire [3:0] n8173_o;
  wire n8175_o;
  wire [3:0] n8176_o;
  wire n8178_o;
  wire n8179_o;
  wire n8180_o;
  wire n8181_o;
  wire n8182_o;
  wire n8183_o;
  wire n8186_o;
  wire n8187_o;
  wire n8190_o;
  wire [6:0] n8191_o;
  wire n8193_o;
  wire n8194_o;
  wire n8195_o;
  wire n8198_o;
  wire n8213_o;
  wire n8215_o;
  wire n8216_o;
  wire n8217_o;
  wire n8218_o;
  wire n8219_o;
  wire n8220_o;
  wire n8221_o;
  wire n8222_o;
  wire n8223_o;
  wire n8224_o;
  wire n8225_o;
  wire n8226_o;
  wire n8227_o;
  wire n8228_o;
  wire n8229_o;
  wire n8230_o;
  wire n8231_o;
  wire n8232_o;
  wire n8233_o;
  wire n8234_o;
  wire n8235_o;
  wire n8236_o;
  wire n8237_o;
  wire n8238_o;
  wire n8239_o;
  wire n8240_o;
  wire n8241_o;
  wire n8244_o;
  wire n8247_o;
  wire n8249_o;
  wire [2:0] n8254_o;
  wire n8258_o;
  wire n8259_o;
  wire n8260_o;
  wire [1:0] n8261_o;
  wire n8264_o;
  wire n8267_o;
  wire n8273_o;
  wire [3:0] n8275_o;
  wire n8283_o;
  wire n8285_o;
  reg n8288_q;
  reg [37:0] n8289_q;
  wire [41:0] n8290_o;
  wire [79:0] n8291_o;
  reg n8292_q;
  wire [89:0] n8293_o;
  wire [7:0] n8294_o;
  reg n8295_q;
  reg [32:0] n8296_q;
  reg [31:0] n8297_q;
  wire [31:0] n8298_o;
  wire [31:0] n8299_o;
  reg [31:0] n8300_q;
  reg n8301_q;
  reg n8302_q;
  reg [39:0] n8303_q;
  reg [3:0] n8304_q;
  wire [218:0] n8305_o;
  reg [6:0] n8306_q;
  reg n8307_q;
  reg [41:0] n8308_q;
  reg [10:0] n8309_q;
  wire [101:0] n8310_o;
  wire [69:0] n8311_o;
  reg [69:0] n8312_q;
  reg [31:0] n8313_q;
  reg n8314_q;
  reg [31:0] n8315_q;
  reg [66:0] n8316_q;
  reg [212:0] n8317_q;
  reg [40:0] n8318_q;
  reg n8319_q;
  wire [497:0] n8320_o;
  reg [31:0] n8322_q;
  reg n8323_q;
  reg [31:0] n8324_q;
  reg [31:0] n8325_q;
  reg n8326_q;
  reg [31:0] n8327_q;
  reg [31:0] n8328_q;
  reg n8329_q;
  reg [31:0] n8330_q;
  reg [31:0] n8331_q;
  reg n8332_q;
  reg [31:0] n8333_q;
  reg [31:0] n8334_q;
  reg n8335_q;
  reg [31:0] n8336_q;
  reg [31:0] n8337_q;
  reg n8338_q;
  reg [31:0] n8339_q;
  reg [31:0] n8340_q;
  reg n8341_q;
  reg [31:0] n8342_q;
  reg [31:0] n8343_q;
  reg n8344_q;
  reg [31:0] n8345_q;
  reg [31:0] n8346_q;
  reg n8347_q;
  reg [31:0] n8348_q;
  reg [31:0] n8349_q;
  reg n8350_q;
  reg [31:0] n8351_q;
  reg [31:0] n8352_q;
  reg n8353_q;
  reg [31:0] n8354_q;
  reg [31:0] n8355_q;
  reg n8356_q;
  reg [31:0] n8357_q;
  reg [31:0] n8358_q;
  reg n8359_q;
  reg [31:0] n8360_q;
  reg [31:0] n8361_q;
  reg n8362_q;
  reg [31:0] n8363_q;
  reg [31:0] n8364_q;
  reg n8365_q;
  reg [31:0] n8366_q;
  reg [31:0] n8367_q;
  reg n8368_q;
  reg [31:0] n8369_q;
  reg [31:0] n8370_q;
  reg n8371_q;
  reg [31:0] n8372_q;
  reg [31:0] n8373_q;
  reg n8374_q;
  reg [31:0] n8375_q;
  reg [31:0] n8376_q;
  reg n8377_q;
  reg [31:0] n8378_q;
  reg [31:0] n8379_q;
  reg n8380_q;
  reg [31:0] n8381_q;
  reg [31:0] n8382_q;
  reg n8383_q;
  reg [31:0] n8384_q;
  reg [31:0] n8385_q;
  reg n8386_q;
  reg [31:0] n8387_q;
  reg [31:0] n8388_q;
  reg n8389_q;
  reg [31:0] n8390_q;
  reg [31:0] n8391_q;
  reg n8392_q;
  reg [31:0] n8393_q;
  reg [31:0] n8394_q;
  reg n8395_q;
  reg [31:0] n8396_q;
  reg [31:0] n8397_q;
  reg n8398_q;
  reg [31:0] n8399_q;
  reg [31:0] n8400_q;
  reg n8401_q;
  reg [31:0] n8402_q;
  reg [31:0] n8403_q;
  reg n8404_q;
  reg [31:0] n8405_q;
  reg [31:0] n8406_q;
  reg n8407_q;
  reg [31:0] n8408_q;
  reg [31:0] n8409_q;
  reg n8410_q;
  reg [31:0] n8411_q;
  reg [31:0] n8412_q;
  reg n8413_q;
  reg [31:0] n8414_q;
  reg [31:0] n8415_q;
  reg n8416_q;
  reg [31:0] n8417_q;
  reg [31:0] n8418_q;
  wire [3231:0] n8419_o;
  wire [1023:0] n8420_o;
  wire [1023:0] n8421_o;
  wire [14:0] n8422_o;
  reg n8423_q;
  reg [1:0] n8424_q;
  wire [8:0] n8425_o;
  wire [69:0] n8426_o;
  reg [31:0] n8427_q;
  wire n8428_o;
  wire n8429_o;
  wire n8430_o;
  wire n8431_o;
  wire n8432_o;
  wire n8433_o;
  wire n8434_o;
  wire n8435_o;
  wire n8436_o;
  wire n8437_o;
  wire n8438_o;
  wire n8439_o;
  wire n8440_o;
  wire n8441_o;
  wire n8442_o;
  wire n8443_o;
  wire n8444_o;
  wire n8445_o;
  wire n8446_o;
  wire n8447_o;
  wire n8448_o;
  wire n8449_o;
  wire n8450_o;
  wire n8451_o;
  wire n8452_o;
  wire n8453_o;
  wire n8454_o;
  wire n8455_o;
  wire n8456_o;
  wire n8457_o;
  wire n8458_o;
  wire n8459_o;
  wire n8460_o;
  wire n8461_o;
  wire n8462_o;
  wire n8463_o;
  wire n8464_o;
  wire n8465_o;
  wire n8466_o;
  wire n8467_o;
  wire n8468_o;
  wire n8469_o;
  wire n8470_o;
  wire n8471_o;
  wire n8472_o;
  wire n8473_o;
  wire n8474_o;
  wire n8475_o;
  wire n8476_o;
  wire n8477_o;
  wire n8478_o;
  wire n8479_o;
  wire n8480_o;
  wire n8481_o;
  wire n8482_o;
  wire n8483_o;
  wire n8484_o;
  wire n8485_o;
  wire n8486_o;
  wire n8487_o;
  wire n8488_o;
  wire n8489_o;
  wire n8490_o;
  wire n8491_o;
  wire n8492_o;
  wire n8493_o;
  wire n8494_o;
  wire n8495_o;
  wire n8496_o;
  wire n8497_o;
  wire n8498_o;
  wire n8499_o;
  wire n8500_o;
  wire n8501_o;
  wire n8502_o;
  wire n8503_o;
  wire n8504_o;
  wire n8505_o;
  wire n8506_o;
  wire n8507_o;
  wire n8508_o;
  wire n8509_o;
  wire n8510_o;
  wire n8511_o;
  wire n8512_o;
  wire n8513_o;
  wire n8514_o;
  wire n8515_o;
  wire n8516_o;
  wire n8517_o;
  wire n8518_o;
  wire n8519_o;
  wire n8520_o;
  wire n8521_o;
  wire n8522_o;
  wire n8523_o;
  wire n8524_o;
  wire n8525_o;
  wire n8526_o;
  wire n8527_o;
  wire n8528_o;
  wire n8529_o;
  wire n8530_o;
  wire n8531_o;
  wire n8532_o;
  wire n8533_o;
  wire n8534_o;
  wire n8535_o;
  wire n8536_o;
  wire n8537_o;
  wire n8538_o;
  wire n8539_o;
  wire n8540_o;
  wire n8541_o;
  wire n8542_o;
  wire n8543_o;
  wire n8544_o;
  wire n8545_o;
  wire n8546_o;
  wire n8547_o;
  wire n8548_o;
  wire n8549_o;
  wire n8550_o;
  wire n8551_o;
  wire n8552_o;
  wire n8553_o;
  wire n8554_o;
  wire n8555_o;
  wire n8556_o;
  wire n8557_o;
  wire n8558_o;
  wire n8559_o;
  wire n8560_o;
  wire n8561_o;
  wire [31:0] n8562_o;
  wire n8563_o;
  wire n8564_o;
  wire n8565_o;
  wire n8566_o;
  wire n8567_o;
  wire n8568_o;
  wire n8569_o;
  wire n8570_o;
  wire n8571_o;
  wire n8572_o;
  wire n8573_o;
  wire n8574_o;
  wire n8575_o;
  wire n8576_o;
  wire n8577_o;
  wire n8578_o;
  wire n8579_o;
  wire n8580_o;
  wire n8581_o;
  wire n8582_o;
  wire n8583_o;
  wire n8584_o;
  wire n8585_o;
  wire n8586_o;
  wire n8587_o;
  wire n8588_o;
  wire n8589_o;
  wire n8590_o;
  wire n8591_o;
  wire n8592_o;
  wire n8593_o;
  wire n8594_o;
  wire n8595_o;
  wire n8596_o;
  wire n8597_o;
  wire n8598_o;
  wire n8599_o;
  wire n8600_o;
  wire n8601_o;
  wire n8602_o;
  wire n8603_o;
  wire n8604_o;
  wire n8605_o;
  wire n8606_o;
  wire n8607_o;
  wire n8608_o;
  wire n8609_o;
  wire n8610_o;
  wire n8611_o;
  wire n8612_o;
  wire n8613_o;
  wire n8614_o;
  wire n8615_o;
  wire n8616_o;
  wire n8617_o;
  wire n8618_o;
  wire n8619_o;
  wire n8620_o;
  wire n8621_o;
  wire n8622_o;
  wire n8623_o;
  wire n8624_o;
  wire n8625_o;
  wire n8626_o;
  wire n8627_o;
  wire n8628_o;
  wire n8629_o;
  wire n8630_o;
  wire n8631_o;
  wire n8632_o;
  wire n8633_o;
  wire n8634_o;
  wire n8635_o;
  wire n8636_o;
  wire n8637_o;
  wire n8638_o;
  wire n8639_o;
  wire n8640_o;
  wire n8641_o;
  wire n8642_o;
  wire n8643_o;
  wire n8644_o;
  wire n8645_o;
  wire n8646_o;
  wire n8647_o;
  wire n8648_o;
  wire n8649_o;
  wire n8650_o;
  wire n8651_o;
  wire n8652_o;
  wire n8653_o;
  wire n8654_o;
  wire n8655_o;
  wire n8656_o;
  wire n8657_o;
  wire n8658_o;
  wire n8659_o;
  wire n8660_o;
  wire n8661_o;
  wire n8662_o;
  wire n8663_o;
  wire n8664_o;
  wire n8665_o;
  wire n8666_o;
  wire n8667_o;
  wire n8668_o;
  wire n8669_o;
  wire n8670_o;
  wire n8671_o;
  wire n8672_o;
  wire n8673_o;
  wire n8674_o;
  wire n8675_o;
  wire n8676_o;
  wire n8677_o;
  wire n8678_o;
  wire n8679_o;
  wire n8680_o;
  wire n8681_o;
  wire n8682_o;
  wire n8683_o;
  wire n8684_o;
  wire n8685_o;
  wire n8686_o;
  wire n8687_o;
  wire n8688_o;
  wire n8689_o;
  wire n8690_o;
  wire n8691_o;
  wire n8692_o;
  wire n8693_o;
  wire n8694_o;
  wire n8695_o;
  wire n8696_o;
  wire [31:0] n8697_o;
  assign ctrl_o_rf_wb_en = n2756_o;
  assign ctrl_o_rf_rs1 = n2757_o;
  assign ctrl_o_rf_rs2 = n2758_o;
  assign ctrl_o_rf_rs3 = n2759_o;
  assign ctrl_o_rf_rd = n2760_o;
  assign ctrl_o_rf_mux = n2761_o;
  assign ctrl_o_rf_zero_we = n2762_o;
  assign ctrl_o_alu_op = n2763_o;
  assign ctrl_o_alu_opa_mux = n2764_o;
  assign ctrl_o_alu_opb_mux = n2765_o;
  assign ctrl_o_alu_unsigned = n2766_o;
  assign ctrl_o_alu_frm = n2767_o;
  assign ctrl_o_alu_cp_trig = n2768_o;
  assign ctrl_o_bus_req = n2769_o;
  assign ctrl_o_bus_mo_we = n2770_o;
  assign ctrl_o_bus_fence = n2771_o;
  assign ctrl_o_bus_fencei = n2772_o;
  assign ctrl_o_bus_priv = n2773_o;
  assign ctrl_o_ir_funct3 = n2774_o;
  assign ctrl_o_ir_funct12 = n2775_o;
  assign ctrl_o_ir_opcode = n2776_o;
  assign ctrl_o_cpu_priv = n2777_o;
  assign ctrl_o_cpu_sleep = n2778_o;
  assign ctrl_o_cpu_trap = n2779_o;
  assign ctrl_o_cpu_debug = n2780_o;
  assign i_bus_addr_o = n2889_o;
  assign i_bus_re_o = n2898_o;
  assign imm_o = n8427_q;
  assign curr_pc_o = n3384_o;
  assign next_pc_o = n3387_o;
  assign csr_rdata_o = n6732_o;
  assign pmp_addr_o = n5681_o;
  assign pmp_ctrl_o = n5680_o;
  assign n2756_o = n8426_o[0];
  assign n2757_o = n8426_o[5:1];
  assign n2758_o = n8426_o[10:6];
  assign n2759_o = n8426_o[15:11];
  assign n2760_o = n8426_o[20:16];
  assign n2761_o = n8426_o[22:21];
  assign n2762_o = n8426_o[23];
  assign n2763_o = n8426_o[26:24];
  assign n2764_o = n8426_o[27];
  assign n2765_o = n8426_o[28];
  assign n2766_o = n8426_o[29];
  assign n2767_o = n8426_o[32:30];
  assign n2768_o = n8426_o[38:33];
  assign n2769_o = n8426_o[39];
  assign n2770_o = n8426_o[40];
  assign n2771_o = n8426_o[41];
  assign n2772_o = n8426_o[42];
  assign n2773_o = n8426_o[43];
  assign n2774_o = n8426_o[46:44];
  assign n2775_o = n8426_o[58:47];
  assign n2776_o = n8426_o[65:59];
  assign n2777_o = n8426_o[66];
  assign n2778_o = n8426_o[67];
  assign n2779_o = n8426_o[68];
  assign n2780_o = n8426_o[69];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:153:10  */
  assign fetch_engine = n8290_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:165:10  */
  assign ipb = n8291_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:178:10  */
  assign issue_engine = n8293_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:191:10  */
  assign decode_aux = n8294_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:224:10  */
  assign execute_engine = n8305_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:246:10  */
  assign trap_ctrl = n8310_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:249:10  */
  assign ctrl_nxt = n8311_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:249:20  */
  assign ctrl = n8312_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:302:10  */
  assign csr = n8320_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:342:10  */
  assign cnt = n8419_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:343:10  */
  assign cnt_lo_rd = n8420_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:344:10  */
  assign cnt_hi_rd = n8421_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:347:10  */
  assign cnt_event = n8422_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:361:10  */
  assign debug_ctrl = n8425_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:364:10  */
  assign illegal_cmd = n4823_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:367:10  */
  assign csr_reg_valid = n4508_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:368:10  */
  assign csr_rw_valid = n4528_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:369:10  */
  assign csr_priv_valid = n4555_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:372:10  */
  assign hw_trigger_fire = n8264_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:375:10  */
  assign imm_opcode = n3268_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:376:10  */
  assign csr_raddr = n6730_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:388:16  */
  assign n2790_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:397:47  */
  assign n2798_o = fetch_engine[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:400:24  */
  assign n2799_o = fetch_engine[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:400:30  */
  assign n2801_o = n2799_o == 2'b00;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:403:46  */
  assign n2803_o = fetch_engine[4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:403:70  */
  assign n2804_o = fetch_engine[38];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:403:54  */
  assign n2805_o = n2803_o | n2804_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:400:7  */
  assign n2806_o = n2801_o ? 1'b0 : n2805_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:407:25  */
  assign n2807_o = fetch_engine[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:411:54  */
  assign n2808_o = execute_engine[116:87];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:411:72  */
  assign n2810_o = {n2808_o, 2'b00};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:412:54  */
  assign n2811_o = execute_engine[86];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:409:9  */
  assign n2814_o = n2807_o == 2'b00;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:418:19  */
  assign n2815_o = ipb[39:38];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:418:24  */
  assign n2817_o = n2815_o == 2'b11;
  assign n2819_o = fetch_engine[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:418:11  */
  assign n2820_o = n2817_o ? 2'b10 : n2819_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:415:9  */
  assign n2822_o = n2807_o == 2'b01;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:424:28  */
  assign n2823_o = fetch_engine[39];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:425:79  */
  assign n2824_o = fetch_engine[37:6];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:425:83  */
  assign n2826_o = n2824_o + 32'b00000000000000000000000000000100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:428:30  */
  assign n2829_o = fetch_engine[4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:428:62  */
  assign n2830_o = fetch_engine[38];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:428:45  */
  assign n2831_o = n2829_o | n2830_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:431:41  */
  assign n2833_o = execute_engine[22:18];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:431:90  */
  assign n2835_o = n2833_o == 5'b11000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:432:41  */
  assign n2836_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:431:121  */
  assign n2837_o = n2835_o & n2836_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:433:40  */
  assign n2838_o = execute_engine[22:18];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:433:89  */
  assign n2840_o = n2838_o == 5'b11011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:432:54  */
  assign n2841_o = n2837_o | n2840_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:434:40  */
  assign n2842_o = execute_engine[22:18];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:434:89  */
  assign n2844_o = n2842_o == 5'b11001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:433:117  */
  assign n2845_o = n2841_o | n2844_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:431:13  */
  assign n2848_o = n2845_o ? 2'b11 : 2'b01;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:428:13  */
  assign n2849_o = n2831_o ? 2'b00 : n2848_o;
  assign n2850_o = {n2826_o, 1'b0};
  assign n2851_o = fetch_engine[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:424:11  */
  assign n2852_o = n2823_o ? n2849_o : n2851_o;
  assign n2853_o = fetch_engine[37:5];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:424:11  */
  assign n2854_o = n2823_o ? n2850_o : n2853_o;
  assign n2855_o = fetch_engine[41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:424:11  */
  assign n2856_o = n2823_o ? 1'b0 : n2855_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:422:9  */
  assign n2858_o = n2807_o == 2'b10;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:443:28  */
  assign n2859_o = fetch_engine[4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:443:60  */
  assign n2860_o = fetch_engine[38];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:443:43  */
  assign n2861_o = n2859_o | n2860_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:443:11  */
  assign n2864_o = n2861_o ? 2'b00 : 2'b01;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:441:9  */
  assign n2866_o = n2807_o == 2'b11;
  assign n2868_o = {n2866_o, n2858_o, n2822_o, n2814_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:407:7  */
  always @*
    case (n2868_o)
      4'b1000: n2869_o = n2864_o;
      4'b0100: n2869_o = n2852_o;
      4'b0010: n2869_o = n2820_o;
      4'b0001: n2869_o = 2'b01;
      default: n2869_o = 2'b00;
    endcase
  assign n2870_o = n2854_o[0];
  assign n2871_o = fetch_engine[5];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:407:7  */
  always @*
    case (n2868_o)
      4'b1000: n2872_o = n2871_o;
      4'b0100: n2872_o = n2870_o;
      4'b0010: n2872_o = n2871_o;
      4'b0001: n2872_o = n2811_o;
      default: n2872_o = n2871_o;
    endcase
  assign n2873_o = n2854_o[32:1];
  assign n2874_o = fetch_engine[37:6];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:407:7  */
  always @*
    case (n2868_o)
      4'b1000: n2875_o = n2874_o;
      4'b0100: n2875_o = n2873_o;
      4'b0010: n2875_o = n2874_o;
      4'b0001: n2875_o = n2810_o;
      default: n2875_o = n2874_o;
    endcase
  assign n2876_o = fetch_engine[41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:407:7  */
  always @*
    case (n2868_o)
      4'b1000: n2877_o = n2876_o;
      4'b0100: n2877_o = n2856_o;
      4'b0010: n2877_o = i_pmp_fault_i;
      4'b0001: n2877_o = n2876_o;
      default: n2877_o = n2876_o;
    endcase
  assign n2878_o = {n2875_o, n2872_o, n2806_o, n2798_o, n2869_o};
  assign n2883_o = {32'b00000000000000000000000000000000, 1'b0, 1'b1, 2'b00, 2'b00};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:458:34  */
  assign n2887_o = fetch_engine[37:8];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:458:52  */
  assign n2889_o = {n2887_o, 2'b00};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:461:40  */
  assign n2891_o = fetch_engine[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:461:46  */
  assign n2893_o = n2891_o == 2'b01;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:461:69  */
  assign n2894_o = ipb[39:38];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:461:74  */
  assign n2896_o = n2894_o == 2'b11;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:461:60  */
  assign n2897_o = n2893_o & n2896_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:461:21  */
  assign n2898_o = n2897_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:464:29  */
  assign n2903_o = 1'b0 ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:468:53  */
  assign n2906_o = i_bus_ack_i | i_bus_err_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:468:28  */
  assign n2907_o = n2906_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:471:48  */
  assign n2909_o = fetch_engine[41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:471:32  */
  assign n2910_o = i_bus_err_i | n2909_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:471:72  */
  assign n2911_o = fetch_engine[40];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:471:57  */
  assign n2912_o = {n2910_o, n2911_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:471:93  */
  assign n2913_o = i_bus_rdata_i[15:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:471:78  */
  assign n2914_o = {n2912_o, n2913_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:472:48  */
  assign n2915_o = fetch_engine[41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:472:32  */
  assign n2916_o = i_bus_err_i | n2915_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:472:72  */
  assign n2917_o = fetch_engine[40];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:472:57  */
  assign n2918_o = {n2916_o, n2917_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:472:93  */
  assign n2919_o = i_bus_rdata_i[31:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:472:78  */
  assign n2920_o = {n2918_o, n2919_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:475:39  */
  assign n2922_o = fetch_engine[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:475:45  */
  assign n2924_o = n2922_o == 2'b10;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:475:77  */
  assign n2925_o = fetch_engine[39];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:475:59  */
  assign n2926_o = n2924_o & n2925_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:476:40  */
  assign n2927_o = fetch_engine[5];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:476:50  */
  assign n2928_o = ~n2927_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:476:57  */
  assign n2930_o = n2928_o | 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:475:89  */
  assign n2931_o = n2926_o & n2930_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:475:20  */
  assign n2932_o = n2931_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:477:39  */
  assign n2935_o = fetch_engine[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:477:45  */
  assign n2937_o = n2935_o == 2'b10;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:477:77  */
  assign n2938_o = fetch_engine[39];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:477:59  */
  assign n2939_o = n2937_o & n2938_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:477:20  */
  assign n2940_o = n2939_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:495:31  */
  assign n2942_o = fetch_engine[4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:498:27  */
  assign n2944_o = ipb[35:18];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:499:24  */
  assign n2945_o = ipb[36];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:500:18  */
  assign prefetch_buffer_n1_prefetch_buffer_inst_n2946 = prefetch_buffer_n1_prefetch_buffer_inst_free_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:502:24  */
  assign n2947_o = ipb[76];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:503:18  */
  assign prefetch_buffer_n1_prefetch_buffer_inst_n2948 = prefetch_buffer_n1_prefetch_buffer_inst_rdata_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:504:18  */
  assign prefetch_buffer_n1_prefetch_buffer_inst_n2949 = prefetch_buffer_n1_prefetch_buffer_inst_avail_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:484:5  */
  neorv32_fifo_2_18_1489f923c4dca729178b3e3233458550d8dddf29 prefetch_buffer_n1_prefetch_buffer_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .clear_i(n2942_o),
    .wdata_i(n2944_o),
    .we_i(n2945_o),
    .re_i(n2947_o),
    .half_o(),
    .free_o(prefetch_buffer_n1_prefetch_buffer_inst_free_o),
    .rdata_o(prefetch_buffer_n1_prefetch_buffer_inst_rdata_o),
    .avail_o(prefetch_buffer_n1_prefetch_buffer_inst_avail_o));
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:495:31  */
  assign n2957_o = fetch_engine[4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:498:27  */
  assign n2959_o = ipb[17:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:499:24  */
  assign n2960_o = ipb[37];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:500:18  */
  assign prefetch_buffer_n2_prefetch_buffer_inst_n2961 = prefetch_buffer_n2_prefetch_buffer_inst_free_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:502:24  */
  assign n2962_o = ipb[77];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:503:18  */
  assign prefetch_buffer_n2_prefetch_buffer_inst_n2963 = prefetch_buffer_n2_prefetch_buffer_inst_rdata_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:504:18  */
  assign prefetch_buffer_n2_prefetch_buffer_inst_n2964 = prefetch_buffer_n2_prefetch_buffer_inst_avail_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:484:5  */
  neorv32_fifo_2_18_1489f923c4dca729178b3e3233458550d8dddf29 prefetch_buffer_n2_prefetch_buffer_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .clear_i(n2957_o),
    .wdata_i(n2959_o),
    .we_i(n2960_o),
    .re_i(n2962_o),
    .half_o(),
    .free_o(prefetch_buffer_n2_prefetch_buffer_inst_free_o),
    .rdata_o(prefetch_buffer_n2_prefetch_buffer_inst_rdata_o),
    .avail_o(prefetch_buffer_n2_prefetch_buffer_inst_avail_o));
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:521:26  */
  assign n2974_o = fetch_engine[4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:522:50  */
  assign n2975_o = execute_engine[86];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:523:31  */
  assign n2976_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:523:37  */
  assign n2978_o = n2976_o == 4'b0001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:524:47  */
  assign n2979_o = issue_engine[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:524:75  */
  assign n2980_o = issue_engine[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:524:58  */
  assign n2981_o = ~n2980_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:524:53  */
  assign n2982_o = n2979_o & n2981_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:524:103  */
  assign n2983_o = issue_engine[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:524:87  */
  assign n2984_o = n2982_o | n2983_o;
  assign n2985_o = issue_engine[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:523:9  */
  assign n2986_o = n2978_o ? n2984_o : n2985_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:521:9  */
  assign n2987_o = n2974_o ? n2975_o : n2986_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:537:24  */
  assign n2995_o = issue_engine[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:537:30  */
  assign n2996_o = ~n2995_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:538:25  */
  assign n2997_o = ipb[59:58];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:538:38  */
  assign n2999_o = n2997_o != 2'b11;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:539:46  */
  assign n3000_o = ipb[78];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:540:46  */
  assign n3001_o = ipb[78];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:541:50  */
  assign n3002_o = issue_engine[51];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:541:71  */
  assign n3003_o = ipb[75:74];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:541:57  */
  assign n3004_o = {n3002_o, n3003_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:541:86  */
  assign n3006_o = {n3004_o, 1'b1};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:541:107  */
  assign n3007_o = issue_engine[50:19];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:541:92  */
  assign n3008_o = {n3006_o, n3007_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:543:54  */
  assign n3009_o = ipb[78];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:543:71  */
  assign n3010_o = ipb[79];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:543:58  */
  assign n3011_o = n3009_o & n3010_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:543:54  */
  assign n3012_o = ipb[78];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:543:71  */
  assign n3013_o = ipb[79];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:543:58  */
  assign n3014_o = n3012_o & n3013_o;
  assign n3015_o = {n3011_o, n3014_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:544:52  */
  assign n3016_o = ipb[57:56];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:544:82  */
  assign n3017_o = ipb[75:74];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:544:67  */
  assign n3018_o = n3016_o | n3017_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:544:37  */
  assign n3020_o = {1'b0, n3018_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:544:98  */
  assign n3022_o = {n3020_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:545:52  */
  assign n3023_o = ipb[55:40];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:545:82  */
  assign n3024_o = ipb[73:58];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:545:68  */
  assign n3025_o = {n3023_o, n3024_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:545:37  */
  assign n3026_o = {n3022_o, n3025_o};
  assign n3027_o = {n3015_o, n3026_o};
  assign n3028_o = {n3001_o, n3008_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:537:7  */
  assign n3029_o = n3076_o ? n3000_o : 1'b0;
  assign n3030_o = n3027_o[36:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:538:9  */
  assign n3031_o = n2999_o ? n3028_o : n3030_o;
  assign n3032_o = n3027_o[37];
  assign n3033_o = n2994_o[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:538:9  */
  assign n3034_o = n2999_o ? n3033_o : n3032_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:549:25  */
  assign n3035_o = ipb[41:40];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:549:38  */
  assign n3037_o = n3035_o != 2'b11;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:550:46  */
  assign n3038_o = ipb[79];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:551:46  */
  assign n3039_o = ipb[79];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:552:50  */
  assign n3040_o = issue_engine[51];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:552:71  */
  assign n3041_o = ipb[57:56];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:552:57  */
  assign n3042_o = {n3040_o, n3041_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:552:86  */
  assign n3044_o = {n3042_o, 1'b1};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:552:107  */
  assign n3045_o = issue_engine[50:19];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:552:92  */
  assign n3046_o = {n3044_o, n3045_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:554:54  */
  assign n3047_o = ipb[78];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:554:71  */
  assign n3048_o = ipb[79];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:554:58  */
  assign n3049_o = n3047_o & n3048_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:554:54  */
  assign n3050_o = ipb[78];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:554:71  */
  assign n3051_o = ipb[79];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:554:58  */
  assign n3052_o = n3050_o & n3051_o;
  assign n3053_o = {n3049_o, n3052_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:555:52  */
  assign n3054_o = ipb[75:74];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:555:82  */
  assign n3055_o = ipb[57:56];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:555:67  */
  assign n3056_o = n3054_o | n3055_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:555:37  */
  assign n3058_o = {1'b0, n3056_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:555:98  */
  assign n3060_o = {n3058_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:556:52  */
  assign n3061_o = ipb[73:58];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:556:82  */
  assign n3062_o = ipb[55:40];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:556:68  */
  assign n3063_o = {n3061_o, n3062_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:556:37  */
  assign n3064_o = {n3060_o, n3063_o};
  assign n3065_o = {n3053_o, n3064_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:549:9  */
  assign n3066_o = n3037_o ? n3038_o : 1'b0;
  assign n3067_o = n3065_o[35:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:549:9  */
  assign n3068_o = n3037_o ? n3046_o : n3067_o;
  assign n3069_o = n3065_o[36];
  assign n3070_o = n2994_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:549:9  */
  assign n3071_o = n3037_o ? n3070_o : n3069_o;
  assign n3072_o = n3065_o[37];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:549:9  */
  assign n3073_o = n3037_o ? n3039_o : n3072_o;
  assign n3074_o = {n3073_o, n3071_o, n3068_o};
  assign n3075_o = {n3034_o, n3031_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:537:7  */
  assign n3076_o = n2996_o & n2999_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:537:7  */
  assign n3077_o = n2996_o ? 1'b0 : n3066_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:537:7  */
  assign n3078_o = n2996_o ? n3075_o : n3074_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:572:44  */
  assign n3081_o = issue_engine[88];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:572:75  */
  assign n3082_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:572:81  */
  assign n3084_o = n3082_o == 4'b0001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:572:55  */
  assign n3085_o = n3081_o & n3084_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:572:20  */
  assign n3086_o = n3085_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:573:44  */
  assign n3089_o = issue_engine[89];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:573:75  */
  assign n3090_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:573:81  */
  assign n3092_o = n3090_o == 4'b0001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:573:55  */
  assign n3093_o = n3089_o & n3092_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:573:20  */
  assign n3094_o = n3093_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:585:36  */
  assign n3096_o = issue_engine[18:3];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:586:23  */
  assign neorv32_cpu_decompressor_inst_true_neorv32_cpu_decompressor_inst_n3097 = neorv32_cpu_decompressor_inst_true_neorv32_cpu_decompressor_inst_ci_illegal_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:587:23  */
  assign neorv32_cpu_decompressor_inst_true_neorv32_cpu_decompressor_inst_n3098 = neorv32_cpu_decompressor_inst_true_neorv32_cpu_decompressor_inst_ci_instr32_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:580:5  */
  neorv32_cpu_decompressor_5ba93c9db0cff93f52b521d7420e43f6eda2784f neorv32_cpu_decompressor_inst_true_neorv32_cpu_decompressor_inst (
    .ci_instr16_i(n3096_o),
    .ci_illegal_o(neorv32_cpu_decompressor_inst_true_neorv32_cpu_decompressor_inst_ci_illegal_o),
    .ci_instr32_o(neorv32_cpu_decompressor_inst_true_neorv32_cpu_decompressor_inst_ci_instr32_o));
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:598:38  */
  assign n3103_o = ipb[73:58];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:598:71  */
  assign n3104_o = issue_engine[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:598:77  */
  assign n3105_o = ~n3104_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:598:52  */
  assign n3106_o = n3105_o ? n3103_o : n3107_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:598:101  */
  assign n3107_o = ipb[55:40];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3110_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3111_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3112_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3113_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3114_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3115_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3116_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3117_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3118_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3119_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3120_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3121_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3122_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3123_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3124_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3125_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3126_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3127_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3128_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3129_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:612:69  */
  assign n3130_o = execute_engine[47];
  assign n3131_o = {n3110_o, n3111_o, n3112_o, n3113_o};
  assign n3132_o = {n3114_o, n3115_o, n3116_o, n3117_o};
  assign n3133_o = {n3118_o, n3119_o, n3120_o, n3121_o};
  assign n3134_o = {n3122_o, n3123_o, n3124_o, n3125_o};
  assign n3135_o = {n3126_o, n3127_o, n3128_o, n3129_o};
  assign n3136_o = {n3131_o, n3132_o, n3133_o, n3134_o};
  assign n3137_o = {n3135_o, n3130_o};
  assign n3138_o = {n3136_o, n3137_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:613:58  */
  assign n3139_o = execute_engine[46:41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:614:58  */
  assign n3140_o = execute_engine[27:23];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:611:9  */
  assign n3142_o = imm_opcode == 7'b0100011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3143_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3144_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3145_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3146_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3147_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3148_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3149_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3150_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3151_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3152_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3153_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3154_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3155_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3156_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3157_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3158_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3159_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3160_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3161_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:616:69  */
  assign n3162_o = execute_engine[47];
  assign n3163_o = {n3143_o, n3144_o, n3145_o, n3146_o};
  assign n3164_o = {n3147_o, n3148_o, n3149_o, n3150_o};
  assign n3165_o = {n3151_o, n3152_o, n3153_o, n3154_o};
  assign n3166_o = {n3155_o, n3156_o, n3157_o, n3158_o};
  assign n3167_o = {n3159_o, n3160_o, n3161_o, n3162_o};
  assign n3168_o = {n3163_o, n3164_o, n3165_o, n3166_o};
  assign n3169_o = {n3168_o, n3167_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:617:58  */
  assign n3170_o = execute_engine[23];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:618:58  */
  assign n3171_o = execute_engine[46:41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:619:58  */
  assign n3172_o = execute_engine[27:24];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:615:9  */
  assign n3175_o = imm_opcode == 7'b1100011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:622:58  */
  assign n3176_o = execute_engine[47:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:621:9  */
  assign n3179_o = imm_opcode == 7'b0110111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:621:27  */
  assign n3181_o = imm_opcode == 7'b0010111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:621:27  */
  assign n3182_o = n3179_o | n3181_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:625:69  */
  assign n3183_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:625:69  */
  assign n3184_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:625:69  */
  assign n3185_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:625:69  */
  assign n3186_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:625:69  */
  assign n3187_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:625:69  */
  assign n3188_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:625:69  */
  assign n3189_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:625:69  */
  assign n3190_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:625:69  */
  assign n3191_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:625:69  */
  assign n3192_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:625:69  */
  assign n3193_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:625:69  */
  assign n3194_o = execute_engine[47];
  assign n3195_o = {n3183_o, n3184_o, n3185_o, n3186_o};
  assign n3196_o = {n3187_o, n3188_o, n3189_o, n3190_o};
  assign n3197_o = {n3191_o, n3192_o, n3193_o, n3194_o};
  assign n3198_o = {n3195_o, n3196_o, n3197_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:626:58  */
  assign n3199_o = execute_engine[35:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:627:58  */
  assign n3200_o = execute_engine[36];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:628:58  */
  assign n3201_o = execute_engine[46:37];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:624:9  */
  assign n3204_o = imm_opcode == 7'b1101111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3205_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3206_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3207_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3208_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3209_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3210_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3211_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3212_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3213_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3214_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3215_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3216_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3217_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3218_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3219_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3220_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3221_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3222_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3223_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3224_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:631:69  */
  assign n3225_o = execute_engine[47];
  assign n3226_o = {n3205_o, n3206_o, n3207_o, n3208_o};
  assign n3227_o = {n3209_o, n3210_o, n3211_o, n3212_o};
  assign n3228_o = {n3213_o, n3214_o, n3215_o, n3216_o};
  assign n3229_o = {n3217_o, n3218_o, n3219_o, n3220_o};
  assign n3230_o = {n3221_o, n3222_o, n3223_o, n3224_o};
  assign n3231_o = {n3226_o, n3227_o, n3228_o, n3229_o};
  assign n3232_o = {n3230_o, n3225_o};
  assign n3233_o = {n3231_o, n3232_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:632:58  */
  assign n3234_o = execute_engine[46:37];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:633:58  */
  assign n3235_o = execute_engine[36];
  assign n3236_o = {n3204_o, n3182_o, n3175_o, n3142_o};
  assign n3237_o = n3140_o[0];
  assign n3238_o = n3177_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:610:7  */
  always @*
    case (n3236_o)
      4'b1000: n3239_o = 1'b0;
      4'b0100: n3239_o = n3238_o;
      4'b0010: n3239_o = 1'b0;
      4'b0001: n3239_o = n3237_o;
      default: n3239_o = n3235_o;
    endcase
  assign n3240_o = n3140_o[4:1];
  assign n3241_o = n3177_o[4:1];
  assign n3242_o = n3201_o[3:0];
  assign n3243_o = n3234_o[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:610:7  */
  always @*
    case (n3236_o)
      4'b1000: n3244_o = n3242_o;
      4'b0100: n3244_o = n3241_o;
      4'b0010: n3244_o = n3172_o;
      4'b0001: n3244_o = n3240_o;
      default: n3244_o = n3243_o;
    endcase
  assign n3245_o = n3177_o[10:5];
  assign n3246_o = n3201_o[9:4];
  assign n3247_o = n3234_o[9:4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:610:7  */
  always @*
    case (n3236_o)
      4'b1000: n3248_o = n3246_o;
      4'b0100: n3248_o = n3245_o;
      4'b0010: n3248_o = n3171_o;
      4'b0001: n3248_o = n3139_o;
      default: n3248_o = n3247_o;
    endcase
  assign n3249_o = n3138_o[0];
  assign n3250_o = n3177_o[11];
  assign n3251_o = n3233_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:610:7  */
  always @*
    case (n3236_o)
      4'b1000: n3252_o = n3200_o;
      4'b0100: n3252_o = n3250_o;
      4'b0010: n3252_o = n3170_o;
      4'b0001: n3252_o = n3249_o;
      default: n3252_o = n3251_o;
    endcase
  assign n3253_o = n3138_o[8:1];
  assign n3254_o = n3169_o[7:0];
  assign n3255_o = n3176_o[7:0];
  assign n3256_o = n3233_o[8:1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:610:7  */
  always @*
    case (n3236_o)
      4'b1000: n3257_o = n3199_o;
      4'b0100: n3257_o = n3255_o;
      4'b0010: n3257_o = n3254_o;
      4'b0001: n3257_o = n3253_o;
      default: n3257_o = n3256_o;
    endcase
  assign n3258_o = n3138_o[20:9];
  assign n3259_o = n3169_o[19:8];
  assign n3260_o = n3176_o[19:8];
  assign n3261_o = n3233_o[20:9];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:610:7  */
  always @*
    case (n3236_o)
      4'b1000: n3262_o = n3198_o;
      4'b0100: n3262_o = n3260_o;
      4'b0010: n3262_o = n3259_o;
      4'b0001: n3262_o = n3258_o;
      default: n3262_o = n3261_o;
    endcase
  assign n3263_o = {n3262_o, n3257_o, n3252_o, n3248_o, n3244_o, n3239_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:639:37  */
  assign n3266_o = execute_engine[22:18];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:639:86  */
  assign n3268_o = {n3266_o, 2'b11};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:646:29  */
  assign n3270_o = execute_engine[30];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:646:50  */
  assign n3271_o = ~n3270_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:647:43  */
  assign n3272_o = cmp_i[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:647:81  */
  assign n3273_o = execute_engine[28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:647:57  */
  assign n3274_o = n3272_o ^ n3273_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:649:43  */
  assign n3275_o = cmp_i[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:649:81  */
  assign n3276_o = execute_engine[28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:649:57  */
  assign n3277_o = n3275_o ^ n3276_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:646:5  */
  assign n3278_o = n3271_o ? n3274_o : n3277_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:658:16  */
  assign n3281_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:673:52  */
  assign n3294_o = execute_engine[7:4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:674:52  */
  assign n3295_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:675:52  */
  assign n3296_o = execute_engine[11:8];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:676:52  */
  assign n3297_o = execute_engine[218];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:677:52  */
  assign n3298_o = execute_engine[79:48];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:678:52  */
  assign n3299_o = execute_engine[81];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:679:52  */
  assign n3300_o = execute_engine[83];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:688:48  */
  assign n3301_o = execute_engine[216];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:692:26  */
  assign n3302_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:692:32  */
  assign n3304_o = n3302_o == 4'b0101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:693:50  */
  assign n3305_o = execute_engine[116:85];
  assign n3306_o = execute_engine[214:183];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:692:7  */
  assign n3307_o = n3304_o ? n3305_o : n3306_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:697:26  */
  assign n3308_o = execute_engine[118];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:698:28  */
  assign n3309_o = execute_engine[117];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:698:39  */
  assign n3310_o = ~n3309_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:699:54  */
  assign n3311_o = execute_engine[150:120];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:699:72  */
  assign n3313_o = {n3311_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:701:41  */
  assign n3314_o = alu_add_i[31:1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:701:59  */
  assign n3316_o = {n3314_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:698:9  */
  assign n3317_o = n3310_o ? n3313_o : n3316_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:706:27  */
  assign n3320_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:713:48  */
  assign n3323_o = csr[191:162];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:713:66  */
  assign n3325_o = {n3323_o, 2'b00};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:707:9  */
  assign n3327_o = n3320_o == 4'b0010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:719:47  */
  assign n3329_o = csr[153:123];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:719:65  */
  assign n3331_o = {n3329_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:715:9  */
  assign n3333_o = n3320_o == 4'b0011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:722:79  */
  assign n3334_o = execute_engine[116:85];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:722:109  */
  assign n3335_o = execute_engine[182:151];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:722:83  */
  assign n3336_o = n3334_o + n3335_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:721:9  */
  assign n3338_o = n3320_o == 4'b0101;
  assign n3339_o = {n3338_o, n3333_o, n3327_o};
  assign n3340_o = execute_engine[150:119];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:706:7  */
  always @*
    case (n3339_o)
      3'b100: n3341_o = n3336_o;
      3'b010: n3341_o = n3331_o;
      3'b001: n3341_o = n3325_o;
      default: n3341_o = n3340_o;
    endcase
  assign n3342_o = {n3298_o, n3296_o, n3295_o};
  assign n3343_o = {n3301_o, n3307_o};
  assign n3361_o = {32'b00000000000000000000000000000000, 4'b0000, 4'b0000};
  assign n3362_o = {1'b0, 32'b00000000000000000000000000000000};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:731:72  */
  assign n3376_o = execute_engine[80];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:731:78  */
  assign n3377_o = ~n3376_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:731:85  */
  assign n3379_o = n3377_o | 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:731:50  */
  assign n3380_o = n3379_o ? 4'b0100 : 4'b0010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:734:33  */
  assign n3382_o = execute_engine[116:86];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:734:51  */
  assign n3384_o = {n3382_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:735:38  */
  assign n3385_o = execute_engine[150:120];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:735:56  */
  assign n3387_o = {n3385_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:743:33  */
  assign n3389_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:743:68  */
  assign n3390_o = trap_ctrl[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:743:47  */
  assign n3391_o = ~n3390_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:743:42  */
  assign n3392_o = n3389_o & n3391_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:744:48  */
  assign n3393_o = execute_engine[35:31];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:745:48  */
  assign n3394_o = execute_engine[40:36];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:746:48  */
  assign n3395_o = execute_engine[47:43];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:747:48  */
  assign n3396_o = execute_engine[27:23];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:748:33  */
  assign n3397_o = ctrl[22:21];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:749:33  */
  assign n3398_o = ctrl[23];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:751:33  */
  assign n3399_o = ctrl[26:24];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:752:33  */
  assign n3400_o = ctrl[27];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:753:33  */
  assign n3401_o = ctrl[28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:754:33  */
  assign n3402_o = ctrl[29];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:755:32  */
  assign n3403_o = csr[322:320];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:756:33  */
  assign n3404_o = ctrl[38:33];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:758:33  */
  assign n3405_o = ctrl[39];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:759:33  */
  assign n3406_o = ctrl[40];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:760:33  */
  assign n3407_o = ctrl[41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:761:33  */
  assign n3408_o = ctrl[42];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:762:13  */
  assign n3409_o = csr[83];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:763:32  */
  assign n3410_o = csr[82];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:765:32  */
  assign n3411_o = csr[121];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:762:5  */
  assign n3412_o = n3409_o ? n3410_o : n3411_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:768:48  */
  assign n3413_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:769:48  */
  assign n3414_o = execute_engine[47:36];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:770:48  */
  assign n3415_o = execute_engine[22:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:772:32  */
  assign n3416_o = csr[121];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:773:43  */
  assign n3417_o = execute_engine[215];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:774:38  */
  assign n3418_o = trap_ctrl[95];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:775:39  */
  assign n3419_o = debug_ctrl[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:851:29  */
  assign n3430_o = execute_engine[47:41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:851:76  */
  assign n3432_o = n3430_o == 7'b0000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:852:106  */
  assign n3433_o = execute_engine[30];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:852:127  */
  assign n3434_o = ~n3433_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:852:81  */
  assign n3436_o = 1'b1 & n3434_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:852:7  */
  assign n3438_o = n3436_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:855:66  */
  assign n3439_o = execute_engine[30];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:855:41  */
  assign n3441_o = 1'b1 & n3439_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:855:7  */
  assign n3443_o = n3441_o ? 1'b1 : 1'b0;
  assign n3444_o = {n3443_o, n3438_o};
  assign n3445_o = {1'b0, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:851:5  */
  assign n3446_o = n3432_o ? n3444_o : n3445_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:867:29  */
  assign n3447_o = execute_engine[35:31];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:867:70  */
  assign n3449_o = n3447_o == 5'b00000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:867:5  */
  assign n3451_o = n3449_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:870:29  */
  assign n3452_o = execute_engine[27:23];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:870:68  */
  assign n3454_o = n3452_o == 5'b00000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:870:5  */
  assign n3456_o = n3454_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:876:35  */
  assign n3458_o = execute_engine[47:36];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:884:51  */
  assign n3460_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:885:51  */
  assign n3461_o = execute_engine[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:886:51  */
  assign n3462_o = execute_engine[80];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:888:51  */
  assign n3464_o = execute_engine[215];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:889:51  */
  assign n3465_o = execute_engine[217];
  assign n3483_o = n3479_o[23];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:914:29  */
  assign n3485_o = execute_engine[20];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:915:52  */
  assign n3486_o = execute_engine[28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:917:52  */
  assign n3487_o = execute_engine[29];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:914:5  */
  assign n3488_o = n3485_o ? n3486_o : n3487_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:25  */
  assign n3491_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:928:57  */
  assign n3493_o = execute_engine[217];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:928:38  */
  assign n3494_o = ~n3493_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:929:55  */
  assign n3495_o = issue_engine[84];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:930:55  */
  assign n3496_o = issue_engine[87];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:932:31  */
  assign n3497_o = issue_engine[88];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:932:64  */
  assign n3498_o = issue_engine[89];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:932:42  */
  assign n3499_o = n3497_o | n3498_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:934:56  */
  assign n3500_o = issue_engine[83:52];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:938:50  */
  assign n3502_o = issue_engine[85];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:938:55  */
  assign n3505_o = n3502_o & 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:939:50  */
  assign n3506_o = issue_engine[86];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:941:30  */
  assign n3507_o = execute_engine[215];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:942:25  */
  assign n3508_o = trap_ctrl[11];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:941:43  */
  assign n3509_o = n3507_o | n3508_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:943:25  */
  assign n3510_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:942:41  */
  assign n3511_o = n3509_o | n3510_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:943:42  */
  assign n3514_o = n3511_o | 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:945:32  */
  assign n3515_o = issue_engine[86];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:944:82  */
  assign n3516_o = n3514_o | n3515_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:941:11  */
  assign n3519_o = n3516_o ? 4'b0010 : 4'b0101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:932:9  */
  assign n3520_o = n3499_o ? n3519_o : n3460_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:932:9  */
  assign n3521_o = n3499_o ? n3500_o : n3461_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:932:9  */
  assign n3522_o = n3499_o ? 1'b0 : n3465_o;
  assign n3523_o = {n3505_o, n3506_o};
  assign n3524_o = {1'b0, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:932:9  */
  assign n3525_o = n3499_o ? n3523_o : n3524_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:924:7  */
  assign n3527_o = n3491_o == 4'b0001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:955:21  */
  assign n3528_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:955:7  */
  assign n3531_o = n3528_o ? 4'b0100 : n3460_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:955:7  */
  assign n3532_o = n3528_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:953:5  */
  assign n3534_o = n3491_o == 4'b0010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:961:7  */
  assign n3538_o = n3491_o == 4'b0011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:967:7  */
  assign n3545_o = n3491_o == 4'b0100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:979:34  */
  assign n3546_o = execute_engine[22:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:984:37  */
  assign n3547_o = execute_engine[21];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:984:60  */
  assign n3548_o = ~n3547_o;
  assign n3550_o = n3479_o[28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:984:13  */
  assign n3551_o = n3548_o ? 1'b1 : n3550_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:989:38  */
  assign n3552_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:991:42  */
  assign n3553_o = execute_engine[21];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:991:97  */
  assign n3554_o = execute_engine[46];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:991:72  */
  assign n3555_o = n3553_o & n3554_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:991:17  */
  assign n3557_o = n3555_o ? 3'b001 : 3'b000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:990:15  */
  assign n3559_o = n3552_o == 3'b000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:996:15  */
  assign n3562_o = n3552_o == 3'b010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:996:33  */
  assign n3564_o = n3552_o == 3'b011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:996:33  */
  assign n3565_o = n3562_o | n3564_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:998:15  */
  assign n3568_o = n3552_o == 3'b100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1000:15  */
  assign n3571_o = n3552_o == 3'b110;
  assign n3573_o = {n3571_o, n3568_o, n3565_o, n3559_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:989:13  */
  always @*
    case (n3573_o)
      4'b1000: n3574_o = 3'b110;
      4'b0100: n3574_o = 3'b101;
      4'b0010: n3574_o = 3'b011;
      4'b0001: n3574_o = n3557_o;
      default: n3574_o = 3'b111;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1007:73  */
  assign n3575_o = execute_engine[21];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1007:48  */
  assign n3577_o = 1'b1 & n3575_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1008:30  */
  assign n3578_o = decode_aux[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1008:61  */
  assign n3579_o = decode_aux[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1008:46  */
  assign n3580_o = n3578_o | n3579_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1007:115  */
  assign n3581_o = n3577_o & n3580_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1008:79  */
  assign n3583_o = n3581_o | 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1025:40  */
  assign n3586_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1025:87  */
  assign n3588_o = n3586_o == 3'b001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1026:40  */
  assign n3589_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1026:87  */
  assign n3591_o = n3589_o == 3'b101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1025:103  */
  assign n3592_o = n3588_o | n3591_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1025:13  */
  assign n3597_o = n3592_o ? 4'b0110 : 4'b0001;
  assign n3598_o = n3479_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1025:13  */
  assign n3599_o = n3592_o ? n3598_o : 1'b1;
  assign n3600_o = n3479_o[33];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1025:13  */
  assign n3601_o = n3592_o ? 1'b1 : n3600_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1007:13  */
  assign n3602_o = n3583_o ? 4'b0110 : n3597_o;
  assign n3603_o = n3479_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1007:13  */
  assign n3604_o = n3583_o ? n3603_o : n3599_o;
  assign n3605_o = n3479_o[33];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1007:13  */
  assign n3606_o = n3583_o ? n3605_o : n3601_o;
  assign n3607_o = n3479_o[34];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1007:13  */
  assign n3608_o = n3583_o ? 1'b1 : n3607_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:981:11  */
  assign n3610_o = n3546_o == 7'b0110011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:981:29  */
  assign n3612_o = n3546_o == 7'b0010011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:981:29  */
  assign n3613_o = n3610_o | n3612_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1040:37  */
  assign n3616_o = execute_engine[21];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1040:13  */
  assign n3618_o = n3616_o ? 3'b100 : 3'b000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1036:11  */
  assign n3622_o = n3546_o == 7'b0110111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1036:29  */
  assign n3624_o = n3546_o == 7'b0010111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1036:29  */
  assign n3625_o = n3622_o | n3624_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1049:11  */
  assign n3630_o = n3546_o == 7'b0000011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1049:30  */
  assign n3632_o = n3546_o == 7'b0100011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1049:30  */
  assign n3633_o = n3630_o | n3632_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1059:37  */
  assign n3635_o = execute_engine[19:18];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1059:88  */
  assign n3637_o = n3635_o == 2'b01;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1059:13  */
  assign n3640_o = n3637_o ? 1'b0 : 1'b1;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1056:11  */
  assign n3643_o = n3546_o == 7'b1100011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1056:32  */
  assign n3645_o = n3546_o == 7'b1101111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1056:32  */
  assign n3646_o = n3643_o | n3645_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1056:47  */
  assign n3648_o = n3546_o == 7'b1100111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1056:47  */
  assign n3649_o = n3646_o | n3648_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1069:37  */
  assign n3650_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1069:84  */
  assign n3652_o = n3650_o == 3'b000;
  assign n3654_o = n3479_o[41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1069:13  */
  assign n3655_o = n3652_o ? 1'b1 : n3654_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1067:11  */
  assign n3661_o = n3546_o == 7'b0001111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1078:11  */
  assign n3664_o = n3546_o == 7'b1010011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1088:11  */
  assign n3667_o = n3546_o == 7'b0001011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1088:31  */
  assign n3669_o = n3546_o == 7'b0101011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1088:31  */
  assign n3670_o = n3667_o | n3669_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1088:48  */
  assign n3672_o = n3546_o == 7'b1011011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1088:48  */
  assign n3673_o = n3670_o | n3672_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1088:65  */
  assign n3675_o = n3546_o == 7'b1111011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1088:65  */
  assign n3676_o = n3673_o | n3675_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1098:11  */
  assign n3680_o = n3546_o == 7'b1110011;
  assign n3682_o = {n3680_o, n3676_o, n3664_o, n3661_o, n3649_o, n3633_o, n3625_o, n3613_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:979:9  */
  always @*
    case (n3682_o)
      8'b10000000: n3683_o = 4'b1000;
      8'b01000000: n3683_o = 4'b0001;
      8'b00100000: n3683_o = 4'b0001;
      8'b00010000: n3683_o = 4'b0100;
      8'b00001000: n3683_o = 4'b0111;
      8'b00000100: n3683_o = 4'b1001;
      8'b00000010: n3683_o = 4'b0001;
      8'b00000001: n3683_o = n3602_o;
      default: n3683_o = 4'b0001;
    endcase
  assign n3684_o = n3479_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:979:9  */
  always @*
    case (n3682_o)
      8'b10000000: n3685_o = n3684_o;
      8'b01000000: n3685_o = n3684_o;
      8'b00100000: n3685_o = n3684_o;
      8'b00010000: n3685_o = n3684_o;
      8'b00001000: n3685_o = n3684_o;
      8'b00000100: n3685_o = n3684_o;
      8'b00000010: n3685_o = 1'b1;
      8'b00000001: n3685_o = n3604_o;
      default: n3685_o = n3684_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:979:9  */
  always @*
    case (n3682_o)
      8'b10000000: n3686_o = 3'b000;
      8'b01000000: n3686_o = 3'b000;
      8'b00100000: n3686_o = 3'b000;
      8'b00010000: n3686_o = 3'b000;
      8'b00001000: n3686_o = 3'b000;
      8'b00000100: n3686_o = 3'b000;
      8'b00000010: n3686_o = n3618_o;
      8'b00000001: n3686_o = n3574_o;
      default: n3686_o = 3'b000;
    endcase
  assign n3687_o = n3479_o[27];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:979:9  */
  always @*
    case (n3682_o)
      8'b10000000: n3688_o = n3687_o;
      8'b01000000: n3688_o = n3687_o;
      8'b00100000: n3688_o = n3687_o;
      8'b00010000: n3688_o = n3687_o;
      8'b00001000: n3688_o = n3640_o;
      8'b00000100: n3688_o = n3687_o;
      8'b00000010: n3688_o = 1'b1;
      8'b00000001: n3688_o = n3687_o;
      default: n3688_o = n3687_o;
    endcase
  assign n3689_o = n3479_o[28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:979:9  */
  always @*
    case (n3682_o)
      8'b10000000: n3690_o = n3689_o;
      8'b01000000: n3690_o = n3689_o;
      8'b00100000: n3690_o = n3689_o;
      8'b00010000: n3690_o = n3689_o;
      8'b00001000: n3690_o = 1'b1;
      8'b00000100: n3690_o = 1'b1;
      8'b00000010: n3690_o = 1'b1;
      8'b00000001: n3690_o = n3551_o;
      default: n3690_o = n3689_o;
    endcase
  assign n3691_o = n3479_o[33];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:979:9  */
  always @*
    case (n3682_o)
      8'b10000000: n3692_o = n3691_o;
      8'b01000000: n3692_o = n3691_o;
      8'b00100000: n3692_o = n3691_o;
      8'b00010000: n3692_o = n3691_o;
      8'b00001000: n3692_o = n3691_o;
      8'b00000100: n3692_o = n3691_o;
      8'b00000010: n3692_o = n3691_o;
      8'b00000001: n3692_o = n3606_o;
      default: n3692_o = n3691_o;
    endcase
  assign n3693_o = n3479_o[34];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:979:9  */
  always @*
    case (n3682_o)
      8'b10000000: n3694_o = n3693_o;
      8'b01000000: n3694_o = n3693_o;
      8'b00100000: n3694_o = n3693_o;
      8'b00010000: n3694_o = n3693_o;
      8'b00001000: n3694_o = n3693_o;
      8'b00000100: n3694_o = n3693_o;
      8'b00000010: n3694_o = n3693_o;
      8'b00000001: n3694_o = n3608_o;
      default: n3694_o = n3693_o;
    endcase
  assign n3695_o = n3479_o[40];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:979:9  */
  always @*
    case (n3682_o)
      8'b10000000: n3696_o = n3695_o;
      8'b01000000: n3696_o = n3695_o;
      8'b00100000: n3696_o = n3695_o;
      8'b00010000: n3696_o = n3695_o;
      8'b00001000: n3696_o = n3695_o;
      8'b00000100: n3696_o = 1'b1;
      8'b00000010: n3696_o = n3695_o;
      8'b00000001: n3696_o = n3695_o;
      default: n3696_o = n3695_o;
    endcase
  assign n3697_o = n3479_o[41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:979:9  */
  always @*
    case (n3682_o)
      8'b10000000: n3698_o = n3697_o;
      8'b01000000: n3698_o = n3697_o;
      8'b00100000: n3698_o = n3697_o;
      8'b00010000: n3698_o = n3655_o;
      8'b00001000: n3698_o = n3697_o;
      8'b00000100: n3698_o = n3697_o;
      8'b00000010: n3698_o = n3697_o;
      8'b00000001: n3698_o = n3697_o;
      default: n3698_o = n3697_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:979:9  */
  always @*
    case (n3682_o)
      8'b10000000: n3699_o = 1'b1;
      8'b01000000: n3699_o = 1'b0;
      8'b00100000: n3699_o = 1'b0;
      8'b00010000: n3699_o = 1'b0;
      8'b00001000: n3699_o = 1'b0;
      8'b00000100: n3699_o = 1'b0;
      8'b00000010: n3699_o = 1'b0;
      8'b00000001: n3699_o = 1'b0;
      default: n3699_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:976:7  */
  assign n3701_o = n3491_o == 4'b0101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1115:55  */
  assign n3703_o = trap_ctrl[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1115:34  */
  assign n3704_o = alu_cp_done_i | n3703_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1115:9  */
  assign n3707_o = n3704_o ? 4'b0001 : n3460_o;
  assign n3708_o = n3479_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1115:9  */
  assign n3709_o = n3704_o ? 1'b1 : n3708_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1111:7  */
  assign n3711_o = n3491_o == 4'b0110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1128:33  */
  assign n3715_o = execute_engine[18];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1128:82  */
  assign n3716_o = execute_engine[84];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1128:63  */
  assign n3717_o = n3715_o | n3716_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1128:9  */
  assign n3721_o = n3717_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1128:9  */
  assign n3722_o = n3717_o ? 4'b0000 : 4'b0001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1135:33  */
  assign n3723_o = execute_engine[18];
  assign n3725_o = n3479_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1135:9  */
  assign n3726_o = n3723_o ? 1'b1 : n3725_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1121:7  */
  assign n3728_o = n3491_o == 4'b0111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1140:7  */
  assign n3734_o = n3491_o == 4'b0000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1153:30  */
  assign n3735_o = trap_ctrl[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1153:47  */
  assign n3736_o = ~n3735_o;
  assign n3738_o = n3479_o[39];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1153:9  */
  assign n3739_o = n3736_o ? 1'b1 : n3738_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1151:7  */
  assign n3742_o = n3491_o == 4'b1001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1163:31  */
  assign n3744_o = trap_ctrl[8];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1163:67  */
  assign n3745_o = trap_ctrl[7];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1163:47  */
  assign n3746_o = n3744_o | n3745_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1164:31  */
  assign n3747_o = trap_ctrl[6];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1163:83  */
  assign n3748_o = n3746_o | n3747_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1164:67  */
  assign n3749_o = trap_ctrl[5];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1164:47  */
  assign n3750_o = n3748_o | n3749_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1165:31  */
  assign n3751_o = trap_ctrl[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1164:83  */
  assign n3752_o = n3750_o | n3751_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1167:29  */
  assign n3754_o = ~bus_d_wait_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1168:35  */
  assign n3755_o = execute_engine[21];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1168:58  */
  assign n3756_o = ~n3755_o;
  assign n3758_o = n3479_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1167:9  */
  assign n3759_o = n3763_o ? 1'b1 : n3758_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1167:9  */
  assign n3761_o = n3754_o ? 4'b0001 : n3460_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1167:9  */
  assign n3763_o = n3754_o & n3756_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1163:9  */
  assign n3764_o = n3752_o ? 4'b0001 : n3761_o;
  assign n3765_o = n3479_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1163:9  */
  assign n3766_o = n3752_o ? n3765_o : n3759_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1159:7  */
  assign n3768_o = n3491_o == 4'b1010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1178:33  */
  assign n3769_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1178:80  */
  assign n3771_o = n3769_o == 3'b000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1179:30  */
  assign n3772_o = trap_ctrl[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1179:47  */
  assign n3773_o = ~n3772_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1178:96  */
  assign n3774_o = n3771_o & n3773_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1181:36  */
  assign n3776_o = execute_engine[47:36];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1182:13  */
  assign n3779_o = n3776_o == 12'b000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1183:13  */
  assign n3782_o = n3776_o == 12'b000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1184:13  */
  assign n3785_o = n3776_o == 12'b001100000010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1185:13  */
  assign n3789_o = n3776_o == 12'b011110110010;
  assign n3791_o = {n3789_o, n3785_o, n3782_o, n3779_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1181:11  */
  always @*
    case (n3791_o)
      4'b1000: n3792_o = 4'b0011;
      4'b0100: n3792_o = 4'b0011;
      4'b0010: n3792_o = 4'b0001;
      4'b0001: n3792_o = 4'b0001;
      default: n3792_o = 4'b0001;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1181:11  */
  always @*
    case (n3791_o)
      4'b1000: n3793_o = n3464_o;
      4'b0100: n3793_o = n3464_o;
      4'b0010: n3793_o = n3464_o;
      4'b0001: n3793_o = n3464_o;
      default: n3793_o = 1'b1;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1181:11  */
  always @*
    case (n3791_o)
      4'b1000: n3794_o = 1'b0;
      4'b0100: n3794_o = 1'b0;
      4'b0010: n3794_o = 1'b0;
      4'b0001: n3794_o = 1'b1;
      default: n3794_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1181:11  */
  always @*
    case (n3791_o)
      4'b1000: n3795_o = 1'b0;
      4'b0100: n3795_o = 1'b0;
      4'b0010: n3795_o = 1'b1;
      4'b0001: n3795_o = 1'b0;
      default: n3795_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1181:11  */
  always @*
    case (n3791_o)
      4'b1000: n3796_o = 1'b1;
      4'b0100: n3796_o = 1'b0;
      4'b0010: n3796_o = 1'b0;
      4'b0001: n3796_o = 1'b0;
      default: n3796_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1190:35  */
  assign n3798_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1190:82  */
  assign n3800_o = n3798_o == 3'b001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1191:35  */
  assign n3801_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1191:82  */
  assign n3803_o = n3801_o == 3'b101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1190:100  */
  assign n3804_o = n3800_o | n3803_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1192:26  */
  assign n3805_o = decode_aux[6];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1192:35  */
  assign n3806_o = ~n3805_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1191:101  */
  assign n3807_o = n3804_o | n3806_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1190:11  */
  assign n3809_o = n3807_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1178:9  */
  assign n3811_o = n3774_o ? n3792_o : 4'b0001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1178:9  */
  assign n3812_o = n3774_o ? n3793_o : n3464_o;
  assign n3813_o = {n3795_o, n3794_o};
  assign n3814_o = {1'b0, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1178:9  */
  assign n3815_o = n3774_o ? n3813_o : n3814_o;
  assign n3816_o = n3479_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1178:9  */
  assign n3817_o = n3774_o ? n3816_o : 1'b1;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1178:9  */
  assign n3818_o = n3774_o ? 1'b0 : n3809_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1178:9  */
  assign n3819_o = n3774_o ? n3796_o : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1175:7  */
  assign n3821_o = n3491_o == 4'b1000;
  assign n3823_o = {n3821_o, n3768_o, n3742_o, n3734_o, n3728_o, n3711_o, n3701_o, n3545_o, n3538_o, n3534_o, n3527_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3824_o = 1'b0;
      11'b01000000000: n3824_o = 1'b0;
      11'b00100000000: n3824_o = 1'b0;
      11'b00010000000: n3824_o = 1'b0;
      11'b00001000000: n3824_o = n3721_o;
      11'b00000100000: n3824_o = 1'b0;
      11'b00000010000: n3824_o = 1'b0;
      11'b00000001000: n3824_o = 1'b1;
      11'b00000000100: n3824_o = 1'b0;
      11'b00000000010: n3824_o = 1'b0;
      11'b00000000001: n3824_o = 1'b0;
      default: n3824_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3825_o = n3811_o;
      11'b01000000000: n3825_o = n3764_o;
      11'b00100000000: n3825_o = 4'b1010;
      11'b00010000000: n3825_o = 4'b0001;
      11'b00001000000: n3825_o = n3722_o;
      11'b00000100000: n3825_o = n3707_o;
      11'b00000010000: n3825_o = n3683_o;
      11'b00000001000: n3825_o = 4'b0000;
      11'b00000000100: n3825_o = 4'b0100;
      11'b00000000010: n3825_o = n3531_o;
      11'b00000000001: n3825_o = n3520_o;
      default: n3825_o = 4'b0001;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3826_o = n3461_o;
      11'b01000000000: n3826_o = n3461_o;
      11'b00100000000: n3826_o = n3461_o;
      11'b00010000000: n3826_o = n3461_o;
      11'b00001000000: n3826_o = n3461_o;
      11'b00000100000: n3826_o = n3461_o;
      11'b00000010000: n3826_o = n3461_o;
      11'b00000001000: n3826_o = n3461_o;
      11'b00000000100: n3826_o = n3461_o;
      11'b00000000010: n3826_o = n3461_o;
      11'b00000000001: n3826_o = n3521_o;
      default: n3826_o = n3461_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3827_o = n3462_o;
      11'b01000000000: n3827_o = n3462_o;
      11'b00100000000: n3827_o = n3462_o;
      11'b00010000000: n3827_o = n3462_o;
      11'b00001000000: n3827_o = n3462_o;
      11'b00000100000: n3827_o = n3462_o;
      11'b00000010000: n3827_o = n3462_o;
      11'b00000001000: n3827_o = n3462_o;
      11'b00000000100: n3827_o = n3462_o;
      11'b00000000010: n3827_o = n3462_o;
      11'b00000000001: n3827_o = n3495_o;
      default: n3827_o = n3462_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3828_o = 1'b0;
      11'b01000000000: n3828_o = 1'b0;
      11'b00100000000: n3828_o = 1'b0;
      11'b00010000000: n3828_o = 1'b0;
      11'b00001000000: n3828_o = 1'b0;
      11'b00000100000: n3828_o = 1'b0;
      11'b00000010000: n3828_o = 1'b0;
      11'b00000001000: n3828_o = 1'b0;
      11'b00000000100: n3828_o = 1'b0;
      11'b00000000010: n3828_o = 1'b0;
      11'b00000000001: n3828_o = n3496_o;
      default: n3828_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3829_o = 1'b0;
      11'b01000000000: n3829_o = 1'b0;
      11'b00100000000: n3829_o = 1'b0;
      11'b00010000000: n3829_o = 1'b0;
      11'b00001000000: n3829_o = 1'b1;
      11'b00000100000: n3829_o = 1'b0;
      11'b00000010000: n3829_o = 1'b0;
      11'b00000001000: n3829_o = 1'b0;
      11'b00000000100: n3829_o = 1'b0;
      11'b00000000010: n3829_o = 1'b0;
      11'b00000000001: n3829_o = 1'b0;
      default: n3829_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3830_o = 1'b0;
      11'b01000000000: n3830_o = 1'b0;
      11'b00100000000: n3830_o = 1'b0;
      11'b00010000000: n3830_o = 1'b0;
      11'b00001000000: n3830_o = 1'b1;
      11'b00000100000: n3830_o = 1'b0;
      11'b00000010000: n3830_o = 1'b0;
      11'b00000001000: n3830_o = 1'b1;
      11'b00000000100: n3830_o = 1'b0;
      11'b00000000010: n3830_o = 1'b0;
      11'b00000000001: n3830_o = n3494_o;
      default: n3830_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3831_o = n3812_o;
      11'b01000000000: n3831_o = n3464_o;
      11'b00100000000: n3831_o = n3464_o;
      11'b00010000000: n3831_o = n3464_o;
      11'b00001000000: n3831_o = n3464_o;
      11'b00000100000: n3831_o = n3464_o;
      11'b00000010000: n3831_o = n3464_o;
      11'b00000001000: n3831_o = 1'b0;
      11'b00000000100: n3831_o = n3464_o;
      11'b00000000010: n3831_o = n3464_o;
      11'b00000000001: n3831_o = n3464_o;
      default: n3831_o = n3464_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3832_o = n3465_o;
      11'b01000000000: n3832_o = n3465_o;
      11'b00100000000: n3832_o = n3465_o;
      11'b00010000000: n3832_o = 1'b1;
      11'b00001000000: n3832_o = n3465_o;
      11'b00000100000: n3832_o = n3465_o;
      11'b00000010000: n3832_o = n3465_o;
      11'b00000001000: n3832_o = n3465_o;
      11'b00000000100: n3832_o = n3465_o;
      11'b00000000010: n3832_o = n3465_o;
      11'b00000000001: n3832_o = n3522_o;
      default: n3832_o = n3465_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3833_o = 1'b0;
      11'b01000000000: n3833_o = 1'b0;
      11'b00100000000: n3833_o = 1'b0;
      11'b00010000000: n3833_o = 1'b0;
      11'b00001000000: n3833_o = 1'b0;
      11'b00000100000: n3833_o = 1'b0;
      11'b00000010000: n3833_o = 1'b0;
      11'b00000001000: n3833_o = 1'b0;
      11'b00000000100: n3833_o = 1'b0;
      11'b00000000010: n3833_o = n3532_o;
      11'b00000000001: n3833_o = 1'b0;
      default: n3833_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3834_o = 1'b0;
      11'b01000000000: n3834_o = 1'b0;
      11'b00100000000: n3834_o = 1'b0;
      11'b00010000000: n3834_o = 1'b0;
      11'b00001000000: n3834_o = 1'b0;
      11'b00000100000: n3834_o = 1'b0;
      11'b00000010000: n3834_o = 1'b0;
      11'b00000001000: n3834_o = 1'b0;
      11'b00000000100: n3834_o = 1'b1;
      11'b00000000010: n3834_o = 1'b0;
      11'b00000000001: n3834_o = 1'b0;
      default: n3834_o = 1'b0;
    endcase
  assign n3835_o = {1'b0, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3836_o = n3835_o;
      11'b01000000000: n3836_o = n3835_o;
      11'b00100000000: n3836_o = n3835_o;
      11'b00010000000: n3836_o = n3835_o;
      11'b00001000000: n3836_o = n3835_o;
      11'b00000100000: n3836_o = n3835_o;
      11'b00000010000: n3836_o = n3835_o;
      11'b00000001000: n3836_o = n3835_o;
      11'b00000000100: n3836_o = n3835_o;
      11'b00000000010: n3836_o = n3835_o;
      11'b00000000001: n3836_o = n3525_o;
      default: n3836_o = n3835_o;
    endcase
  assign n3837_o = {1'b0, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3838_o = n3815_o;
      11'b01000000000: n3838_o = n3837_o;
      11'b00100000000: n3838_o = n3837_o;
      11'b00010000000: n3838_o = n3837_o;
      11'b00001000000: n3838_o = n3837_o;
      11'b00000100000: n3838_o = n3837_o;
      11'b00000010000: n3838_o = n3837_o;
      11'b00000001000: n3838_o = n3837_o;
      11'b00000000100: n3838_o = n3837_o;
      11'b00000000010: n3838_o = n3837_o;
      11'b00000000001: n3838_o = n3837_o;
      default: n3838_o = n3837_o;
    endcase
  assign n3839_o = n3479_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3840_o = n3817_o;
      11'b01000000000: n3840_o = n3766_o;
      11'b00100000000: n3840_o = n3839_o;
      11'b00010000000: n3840_o = n3839_o;
      11'b00001000000: n3840_o = n3726_o;
      11'b00000100000: n3840_o = n3709_o;
      11'b00000010000: n3840_o = n3685_o;
      11'b00000001000: n3840_o = n3839_o;
      11'b00000000100: n3840_o = n3839_o;
      11'b00000000010: n3840_o = n3839_o;
      11'b00000000001: n3840_o = n3839_o;
      default: n3840_o = n3839_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3841_o = 2'b10;
      11'b01000000000: n3841_o = 2'b01;
      11'b00100000000: n3841_o = 2'b00;
      11'b00010000000: n3841_o = 2'b10;
      11'b00001000000: n3841_o = 2'b11;
      11'b00000100000: n3841_o = 2'b00;
      11'b00000010000: n3841_o = 2'b00;
      11'b00000001000: n3841_o = 2'b00;
      11'b00000000100: n3841_o = 2'b00;
      11'b00000000010: n3841_o = 2'b00;
      11'b00000000001: n3841_o = 2'b00;
      default: n3841_o = 2'b00;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3842_o = n3483_o;
      11'b01000000000: n3842_o = n3483_o;
      11'b00100000000: n3842_o = n3483_o;
      11'b00010000000: n3842_o = 1'b1;
      11'b00001000000: n3842_o = n3483_o;
      11'b00000100000: n3842_o = n3483_o;
      11'b00000010000: n3842_o = n3483_o;
      11'b00000001000: n3842_o = n3483_o;
      11'b00000000100: n3842_o = n3483_o;
      11'b00000000010: n3842_o = n3483_o;
      11'b00000000001: n3842_o = n3483_o;
      default: n3842_o = n3483_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3843_o = 3'b000;
      11'b01000000000: n3843_o = 3'b000;
      11'b00100000000: n3843_o = 3'b000;
      11'b00010000000: n3843_o = 3'b000;
      11'b00001000000: n3843_o = 3'b000;
      11'b00000100000: n3843_o = 3'b010;
      11'b00000010000: n3843_o = n3686_o;
      11'b00000001000: n3843_o = 3'b000;
      11'b00000000100: n3843_o = 3'b000;
      11'b00000000010: n3843_o = 3'b000;
      11'b00000000001: n3843_o = 3'b000;
      default: n3843_o = 3'b000;
    endcase
  assign n3844_o = n3479_o[27];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3845_o = n3844_o;
      11'b01000000000: n3845_o = n3844_o;
      11'b00100000000: n3845_o = n3844_o;
      11'b00010000000: n3845_o = n3844_o;
      11'b00001000000: n3845_o = n3844_o;
      11'b00000100000: n3845_o = n3844_o;
      11'b00000010000: n3845_o = n3688_o;
      11'b00000001000: n3845_o = n3844_o;
      11'b00000000100: n3845_o = n3844_o;
      11'b00000000010: n3845_o = n3844_o;
      11'b00000000001: n3845_o = n3844_o;
      default: n3845_o = n3844_o;
    endcase
  assign n3846_o = n3479_o[28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3847_o = n3846_o;
      11'b01000000000: n3847_o = n3846_o;
      11'b00100000000: n3847_o = n3846_o;
      11'b00010000000: n3847_o = n3846_o;
      11'b00001000000: n3847_o = n3846_o;
      11'b00000100000: n3847_o = n3846_o;
      11'b00000010000: n3847_o = n3690_o;
      11'b00000001000: n3847_o = n3846_o;
      11'b00000000100: n3847_o = n3846_o;
      11'b00000000010: n3847_o = n3846_o;
      11'b00000000001: n3847_o = n3846_o;
      default: n3847_o = n3846_o;
    endcase
  assign n3848_o = n3479_o[33];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3849_o = n3848_o;
      11'b01000000000: n3849_o = n3848_o;
      11'b00100000000: n3849_o = n3848_o;
      11'b00010000000: n3849_o = n3848_o;
      11'b00001000000: n3849_o = n3848_o;
      11'b00000100000: n3849_o = n3848_o;
      11'b00000010000: n3849_o = n3692_o;
      11'b00000001000: n3849_o = n3848_o;
      11'b00000000100: n3849_o = n3848_o;
      11'b00000000010: n3849_o = n3848_o;
      11'b00000000001: n3849_o = n3848_o;
      default: n3849_o = n3848_o;
    endcase
  assign n3850_o = n3479_o[34];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3851_o = n3850_o;
      11'b01000000000: n3851_o = n3850_o;
      11'b00100000000: n3851_o = n3850_o;
      11'b00010000000: n3851_o = n3850_o;
      11'b00001000000: n3851_o = n3850_o;
      11'b00000100000: n3851_o = n3850_o;
      11'b00000010000: n3851_o = n3694_o;
      11'b00000001000: n3851_o = n3850_o;
      11'b00000000100: n3851_o = n3850_o;
      11'b00000000010: n3851_o = n3850_o;
      11'b00000000001: n3851_o = n3850_o;
      default: n3851_o = n3850_o;
    endcase
  assign n3852_o = n3479_o[39];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3853_o = n3852_o;
      11'b01000000000: n3853_o = n3852_o;
      11'b00100000000: n3853_o = n3739_o;
      11'b00010000000: n3853_o = n3852_o;
      11'b00001000000: n3853_o = n3852_o;
      11'b00000100000: n3853_o = n3852_o;
      11'b00000010000: n3853_o = n3852_o;
      11'b00000001000: n3853_o = n3852_o;
      11'b00000000100: n3853_o = n3852_o;
      11'b00000000010: n3853_o = n3852_o;
      11'b00000000001: n3853_o = n3852_o;
      default: n3853_o = n3852_o;
    endcase
  assign n3854_o = n3479_o[40];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3855_o = n3854_o;
      11'b01000000000: n3855_o = n3854_o;
      11'b00100000000: n3855_o = n3854_o;
      11'b00010000000: n3855_o = n3854_o;
      11'b00001000000: n3855_o = n3854_o;
      11'b00000100000: n3855_o = n3854_o;
      11'b00000010000: n3855_o = n3696_o;
      11'b00000001000: n3855_o = n3854_o;
      11'b00000000100: n3855_o = n3854_o;
      11'b00000000010: n3855_o = n3854_o;
      11'b00000000001: n3855_o = n3854_o;
      default: n3855_o = n3854_o;
    endcase
  assign n3856_o = n3479_o[41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3857_o = n3856_o;
      11'b01000000000: n3857_o = n3856_o;
      11'b00100000000: n3857_o = n3856_o;
      11'b00010000000: n3857_o = n3856_o;
      11'b00001000000: n3857_o = n3856_o;
      11'b00000100000: n3857_o = n3856_o;
      11'b00000010000: n3857_o = n3698_o;
      11'b00000001000: n3857_o = n3856_o;
      11'b00000000100: n3857_o = n3856_o;
      11'b00000000010: n3857_o = n3856_o;
      11'b00000000001: n3857_o = n3856_o;
      default: n3857_o = n3856_o;
    endcase
  assign n3858_o = n3479_o[20:1];
  assign n3861_o = n3479_o[32:30];
  assign n3864_o = n3479_o[38:35];
  assign n3866_o = n3479_o[69:42];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3867_o = n3818_o;
      11'b01000000000: n3867_o = 1'b0;
      11'b00100000000: n3867_o = 1'b0;
      11'b00010000000: n3867_o = 1'b0;
      11'b00001000000: n3867_o = 1'b0;
      11'b00000100000: n3867_o = 1'b0;
      11'b00000010000: n3867_o = 1'b0;
      11'b00000001000: n3867_o = 1'b0;
      11'b00000000100: n3867_o = 1'b0;
      11'b00000000010: n3867_o = 1'b0;
      11'b00000000001: n3867_o = 1'b0;
      default: n3867_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3868_o = 1'b0;
      11'b01000000000: n3868_o = 1'b0;
      11'b00100000000: n3868_o = 1'b0;
      11'b00010000000: n3868_o = 1'b0;
      11'b00001000000: n3868_o = 1'b0;
      11'b00000100000: n3868_o = 1'b0;
      11'b00000010000: n3868_o = n3699_o;
      11'b00000001000: n3868_o = 1'b0;
      11'b00000000100: n3868_o = 1'b0;
      11'b00000000010: n3868_o = 1'b0;
      11'b00000000001: n3868_o = 1'b0;
      default: n3868_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:922:5  */
  always @*
    case (n3823_o)
      11'b10000000000: n3869_o = n3819_o;
      11'b01000000000: n3869_o = 1'b0;
      11'b00100000000: n3869_o = 1'b0;
      11'b00010000000: n3869_o = 1'b0;
      11'b00001000000: n3869_o = 1'b0;
      11'b00000100000: n3869_o = 1'b0;
      11'b00000010000: n3869_o = 1'b0;
      11'b00000001000: n3869_o = 1'b0;
      11'b00000000100: n3869_o = 1'b0;
      11'b00000000010: n3869_o = 1'b0;
      11'b00000000001: n3869_o = 1'b0;
      default: n3869_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1216:14  */
  assign n3872_o = csr[11:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1219:7  */
  assign n3875_o = n3872_o == 12'b000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1219:25  */
  assign n3877_o = n3872_o == 12'b000000000010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1219:25  */
  assign n3878_o = n3875_o | n3877_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1219:37  */
  assign n3880_o = n3872_o == 12'b000000000011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1219:37  */
  assign n3881_o = n3878_o | n3880_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1223:7  */
  assign n3883_o = n3872_o == 12'b001100000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1223:26  */
  assign n3885_o = n3872_o == 12'b001100010000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1223:26  */
  assign n3886_o = n3883_o | n3885_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1223:43  */
  assign n3888_o = n3872_o == 12'b001100000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1223:43  */
  assign n3889_o = n3886_o | n3888_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1223:56  */
  assign n3891_o = n3872_o == 12'b001100000100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1223:56  */
  assign n3892_o = n3889_o | n3891_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1223:68  */
  assign n3894_o = n3872_o == 12'b001100000101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1223:68  */
  assign n3895_o = n3892_o | n3894_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1223:82  */
  assign n3897_o = n3872_o == 12'b001101000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1223:82  */
  assign n3898_o = n3895_o | n3897_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1223:99  */
  assign n3900_o = n3872_o == 12'b001101000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1223:99  */
  assign n3901_o = n3898_o | n3900_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1223:112  */
  assign n3903_o = n3872_o == 12'b001101000010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1223:112  */
  assign n3904_o = n3901_o | n3903_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1224:25  */
  assign n3906_o = n3872_o == 12'b001101000100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1224:25  */
  assign n3907_o = n3904_o | n3906_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1224:37  */
  assign n3909_o = n3872_o == 12'b001101000011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1224:37  */
  assign n3910_o = n3907_o | n3909_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1224:51  */
  assign n3912_o = n3872_o == 12'b001100100000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1224:51  */
  assign n3913_o = n3910_o | n3912_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1224:73  */
  assign n3915_o = n3872_o == 12'b001100000110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1224:73  */
  assign n3916_o = n3913_o | n3915_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1224:92  */
  assign n3918_o = n3872_o == 12'b001100001010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1224:92  */
  assign n3919_o = n3916_o | n3918_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1224:108  */
  assign n3921_o = n3872_o == 12'b001100011010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1224:108  */
  assign n3922_o = n3919_o | n3921_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1224:125  */
  assign n3924_o = n3872_o == 12'b111100010001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1224:125  */
  assign n3925_o = n3922_o | n3924_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1225:28  */
  assign n3927_o = n3872_o == 12'b111100010010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1225:28  */
  assign n3928_o = n3925_o | n3927_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1225:44  */
  assign n3930_o = n3872_o == 12'b111100010011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1225:44  */
  assign n3931_o = n3928_o | n3930_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1225:59  */
  assign n3933_o = n3872_o == 12'b111100010100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1225:59  */
  assign n3934_o = n3931_o | n3933_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1225:75  */
  assign n3936_o = n3872_o == 12'b111100010101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1225:75  */
  assign n3937_o = n3934_o | n3936_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1225:94  */
  assign n3939_o = n3872_o == 12'b111111000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1225:94  */
  assign n3940_o = n3937_o | n3939_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1229:7  */
  assign n3943_o = n3872_o == 12'b001110110000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1229:27  */
  assign n3945_o = n3872_o == 12'b001110110001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1229:27  */
  assign n3946_o = n3943_o | n3945_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1229:44  */
  assign n3948_o = n3872_o == 12'b001110110010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1229:44  */
  assign n3949_o = n3946_o | n3948_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1229:62  */
  assign n3951_o = n3872_o == 12'b001110110011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1229:62  */
  assign n3952_o = n3949_o | n3951_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1229:80  */
  assign n3954_o = n3872_o == 12'b001110110100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1229:80  */
  assign n3955_o = n3952_o | n3954_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1229:98  */
  assign n3957_o = n3872_o == 12'b001110110101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1229:98  */
  assign n3958_o = n3955_o | n3957_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1229:116  */
  assign n3960_o = n3872_o == 12'b001110110110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1229:116  */
  assign n3961_o = n3958_o | n3960_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1229:134  */
  assign n3963_o = n3872_o == 12'b001110110111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1229:134  */
  assign n3964_o = n3961_o | n3963_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1229:152  */
  assign n3966_o = n3872_o == 12'b001110111000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1229:152  */
  assign n3967_o = n3964_o | n3966_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1230:27  */
  assign n3969_o = n3872_o == 12'b001110111001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1230:27  */
  assign n3970_o = n3967_o | n3969_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1230:44  */
  assign n3972_o = n3872_o == 12'b001110111010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1230:44  */
  assign n3973_o = n3970_o | n3972_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1230:62  */
  assign n3975_o = n3872_o == 12'b001110111011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1230:62  */
  assign n3976_o = n3973_o | n3975_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1230:80  */
  assign n3978_o = n3872_o == 12'b001110111100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1230:80  */
  assign n3979_o = n3976_o | n3978_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1230:98  */
  assign n3981_o = n3872_o == 12'b001110111101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1230:98  */
  assign n3982_o = n3979_o | n3981_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1230:116  */
  assign n3984_o = n3872_o == 12'b001110111110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1230:116  */
  assign n3985_o = n3982_o | n3984_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1230:134  */
  assign n3987_o = n3872_o == 12'b001110111111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1230:134  */
  assign n3988_o = n3985_o | n3987_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1230:152  */
  assign n3990_o = n3872_o == 12'b001110100000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1230:152  */
  assign n3991_o = n3988_o | n3990_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1231:27  */
  assign n3993_o = n3872_o == 12'b001110100001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1231:27  */
  assign n3994_o = n3991_o | n3993_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1231:44  */
  assign n3996_o = n3872_o == 12'b001110100010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1231:44  */
  assign n3997_o = n3994_o | n3996_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1231:62  */
  assign n3999_o = n3872_o == 12'b001110100011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1231:62  */
  assign n4000_o = n3997_o | n3999_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1235:7  */
  assign n4003_o = n3872_o == 12'b110000000011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1235:33  */
  assign n4005_o = n3872_o == 12'b110000000100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1235:33  */
  assign n4006_o = n4003_o | n4005_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1235:56  */
  assign n4008_o = n3872_o == 12'b110000000101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1235:56  */
  assign n4009_o = n4006_o | n4008_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1235:79  */
  assign n4011_o = n3872_o == 12'b110000000110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1235:79  */
  assign n4012_o = n4009_o | n4011_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1235:102  */
  assign n4014_o = n3872_o == 12'b110000000111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1235:102  */
  assign n4015_o = n4012_o | n4014_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1235:125  */
  assign n4017_o = n3872_o == 12'b110000001000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1235:125  */
  assign n4018_o = n4015_o | n4017_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1235:148  */
  assign n4020_o = n3872_o == 12'b110000001001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1235:148  */
  assign n4021_o = n4018_o | n4020_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1236:33  */
  assign n4023_o = n3872_o == 12'b110000001010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1236:33  */
  assign n4024_o = n4021_o | n4023_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1236:56  */
  assign n4026_o = n3872_o == 12'b110000001011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1236:56  */
  assign n4027_o = n4024_o | n4026_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1236:79  */
  assign n4029_o = n3872_o == 12'b110000001100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1236:79  */
  assign n4030_o = n4027_o | n4029_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1236:102  */
  assign n4032_o = n3872_o == 12'b110000001101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1236:102  */
  assign n4033_o = n4030_o | n4032_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1236:125  */
  assign n4035_o = n3872_o == 12'b110000001110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1236:125  */
  assign n4036_o = n4033_o | n4035_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1236:148  */
  assign n4038_o = n3872_o == 12'b110000001111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1236:148  */
  assign n4039_o = n4036_o | n4038_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1237:33  */
  assign n4041_o = n3872_o == 12'b110000010000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1237:33  */
  assign n4042_o = n4039_o | n4041_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1237:56  */
  assign n4044_o = n3872_o == 12'b110000010001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1237:56  */
  assign n4045_o = n4042_o | n4044_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1237:79  */
  assign n4047_o = n3872_o == 12'b110000010010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1237:79  */
  assign n4048_o = n4045_o | n4047_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1237:102  */
  assign n4050_o = n3872_o == 12'b110000010011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1237:102  */
  assign n4051_o = n4048_o | n4050_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1237:125  */
  assign n4053_o = n3872_o == 12'b110000010100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1237:125  */
  assign n4054_o = n4051_o | n4053_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1237:148  */
  assign n4056_o = n3872_o == 12'b110000010101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1237:148  */
  assign n4057_o = n4054_o | n4056_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1238:33  */
  assign n4059_o = n3872_o == 12'b110000010110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1238:33  */
  assign n4060_o = n4057_o | n4059_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1238:56  */
  assign n4062_o = n3872_o == 12'b110000010111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1238:56  */
  assign n4063_o = n4060_o | n4062_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1238:79  */
  assign n4065_o = n3872_o == 12'b110000011000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1238:79  */
  assign n4066_o = n4063_o | n4065_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1238:102  */
  assign n4068_o = n3872_o == 12'b110000011001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1238:102  */
  assign n4069_o = n4066_o | n4068_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1238:125  */
  assign n4071_o = n3872_o == 12'b110000011010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1238:125  */
  assign n4072_o = n4069_o | n4071_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1238:148  */
  assign n4074_o = n3872_o == 12'b110000011011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1238:148  */
  assign n4075_o = n4072_o | n4074_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1239:33  */
  assign n4077_o = n3872_o == 12'b110000011100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1239:33  */
  assign n4078_o = n4075_o | n4077_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1239:56  */
  assign n4080_o = n3872_o == 12'b110000011101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1239:56  */
  assign n4081_o = n4078_o | n4080_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1239:79  */
  assign n4083_o = n3872_o == 12'b110000011110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1239:79  */
  assign n4084_o = n4081_o | n4083_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1239:102  */
  assign n4086_o = n3872_o == 12'b110000011111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1239:102  */
  assign n4087_o = n4084_o | n4086_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1239:125  */
  assign n4089_o = n3872_o == 12'b110010000011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1239:125  */
  assign n4090_o = n4087_o | n4089_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1240:33  */
  assign n4092_o = n3872_o == 12'b110010000100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1240:33  */
  assign n4093_o = n4090_o | n4092_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1240:56  */
  assign n4095_o = n3872_o == 12'b110010000101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1240:56  */
  assign n4096_o = n4093_o | n4095_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1240:79  */
  assign n4098_o = n3872_o == 12'b110010000110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1240:79  */
  assign n4099_o = n4096_o | n4098_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1240:102  */
  assign n4101_o = n3872_o == 12'b110010000111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1240:102  */
  assign n4102_o = n4099_o | n4101_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1240:125  */
  assign n4104_o = n3872_o == 12'b110010001000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1240:125  */
  assign n4105_o = n4102_o | n4104_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1240:148  */
  assign n4107_o = n3872_o == 12'b110010001001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1240:148  */
  assign n4108_o = n4105_o | n4107_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1241:33  */
  assign n4110_o = n3872_o == 12'b110010001010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1241:33  */
  assign n4111_o = n4108_o | n4110_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1241:56  */
  assign n4113_o = n3872_o == 12'b110010001011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1241:56  */
  assign n4114_o = n4111_o | n4113_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1241:79  */
  assign n4116_o = n3872_o == 12'b110010001100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1241:79  */
  assign n4117_o = n4114_o | n4116_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1241:102  */
  assign n4119_o = n3872_o == 12'b110010001101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1241:102  */
  assign n4120_o = n4117_o | n4119_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1241:125  */
  assign n4122_o = n3872_o == 12'b110010001110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1241:125  */
  assign n4123_o = n4120_o | n4122_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1241:148  */
  assign n4125_o = n3872_o == 12'b110010001111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1241:148  */
  assign n4126_o = n4123_o | n4125_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1242:33  */
  assign n4128_o = n3872_o == 12'b110010010000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1242:33  */
  assign n4129_o = n4126_o | n4128_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1242:56  */
  assign n4131_o = n3872_o == 12'b110010010001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1242:56  */
  assign n4132_o = n4129_o | n4131_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1242:79  */
  assign n4134_o = n3872_o == 12'b110010010010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1242:79  */
  assign n4135_o = n4132_o | n4134_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1242:102  */
  assign n4137_o = n3872_o == 12'b110010010011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1242:102  */
  assign n4138_o = n4135_o | n4137_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1242:125  */
  assign n4140_o = n3872_o == 12'b110010010100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1242:125  */
  assign n4141_o = n4138_o | n4140_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1242:148  */
  assign n4143_o = n3872_o == 12'b110010010101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1242:148  */
  assign n4144_o = n4141_o | n4143_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1243:33  */
  assign n4146_o = n3872_o == 12'b110010010110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1243:33  */
  assign n4147_o = n4144_o | n4146_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1243:56  */
  assign n4149_o = n3872_o == 12'b110010010111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1243:56  */
  assign n4150_o = n4147_o | n4149_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1243:79  */
  assign n4152_o = n3872_o == 12'b110010011000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1243:79  */
  assign n4153_o = n4150_o | n4152_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1243:102  */
  assign n4155_o = n3872_o == 12'b110010011001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1243:102  */
  assign n4156_o = n4153_o | n4155_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1243:125  */
  assign n4158_o = n3872_o == 12'b110010011010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1243:125  */
  assign n4159_o = n4156_o | n4158_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1243:148  */
  assign n4161_o = n3872_o == 12'b110010011011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1243:148  */
  assign n4162_o = n4159_o | n4161_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1244:33  */
  assign n4164_o = n3872_o == 12'b110010011100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1244:33  */
  assign n4165_o = n4162_o | n4164_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1244:56  */
  assign n4167_o = n3872_o == 12'b110010011101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1244:56  */
  assign n4168_o = n4165_o | n4167_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1244:79  */
  assign n4170_o = n3872_o == 12'b110010011110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1244:79  */
  assign n4171_o = n4168_o | n4170_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1244:102  */
  assign n4173_o = n3872_o == 12'b110010011111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1244:102  */
  assign n4174_o = n4171_o | n4173_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1244:125  */
  assign n4176_o = n3872_o == 12'b101100000011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1244:125  */
  assign n4177_o = n4174_o | n4176_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1245:33  */
  assign n4179_o = n3872_o == 12'b101100000100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1245:33  */
  assign n4180_o = n4177_o | n4179_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1245:56  */
  assign n4182_o = n3872_o == 12'b101100000101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1245:56  */
  assign n4183_o = n4180_o | n4182_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1245:79  */
  assign n4185_o = n3872_o == 12'b101100000110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1245:79  */
  assign n4186_o = n4183_o | n4185_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1245:102  */
  assign n4188_o = n3872_o == 12'b101100000111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1245:102  */
  assign n4189_o = n4186_o | n4188_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1245:125  */
  assign n4191_o = n3872_o == 12'b101100001000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1245:125  */
  assign n4192_o = n4189_o | n4191_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1245:148  */
  assign n4194_o = n3872_o == 12'b101100001001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1245:148  */
  assign n4195_o = n4192_o | n4194_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1246:33  */
  assign n4197_o = n3872_o == 12'b101100001010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1246:33  */
  assign n4198_o = n4195_o | n4197_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1246:56  */
  assign n4200_o = n3872_o == 12'b101100001011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1246:56  */
  assign n4201_o = n4198_o | n4200_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1246:79  */
  assign n4203_o = n3872_o == 12'b101100001100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1246:79  */
  assign n4204_o = n4201_o | n4203_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1246:102  */
  assign n4206_o = n3872_o == 12'b101100001101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1246:102  */
  assign n4207_o = n4204_o | n4206_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1246:125  */
  assign n4209_o = n3872_o == 12'b101100001110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1246:125  */
  assign n4210_o = n4207_o | n4209_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1246:148  */
  assign n4212_o = n3872_o == 12'b101100001111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1246:148  */
  assign n4213_o = n4210_o | n4212_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1247:33  */
  assign n4215_o = n3872_o == 12'b101100010000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1247:33  */
  assign n4216_o = n4213_o | n4215_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1247:56  */
  assign n4218_o = n3872_o == 12'b101100010001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1247:56  */
  assign n4219_o = n4216_o | n4218_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1247:79  */
  assign n4221_o = n3872_o == 12'b101100010010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1247:79  */
  assign n4222_o = n4219_o | n4221_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1247:102  */
  assign n4224_o = n3872_o == 12'b101100010011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1247:102  */
  assign n4225_o = n4222_o | n4224_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1247:125  */
  assign n4227_o = n3872_o == 12'b101100010100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1247:125  */
  assign n4228_o = n4225_o | n4227_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1247:148  */
  assign n4230_o = n3872_o == 12'b101100010101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1247:148  */
  assign n4231_o = n4228_o | n4230_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1248:33  */
  assign n4233_o = n3872_o == 12'b101100010110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1248:33  */
  assign n4234_o = n4231_o | n4233_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1248:56  */
  assign n4236_o = n3872_o == 12'b101100010111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1248:56  */
  assign n4237_o = n4234_o | n4236_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1248:79  */
  assign n4239_o = n3872_o == 12'b101100011000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1248:79  */
  assign n4240_o = n4237_o | n4239_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1248:102  */
  assign n4242_o = n3872_o == 12'b101100011001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1248:102  */
  assign n4243_o = n4240_o | n4242_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1248:125  */
  assign n4245_o = n3872_o == 12'b101100011010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1248:125  */
  assign n4246_o = n4243_o | n4245_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1248:148  */
  assign n4248_o = n3872_o == 12'b101100011011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1248:148  */
  assign n4249_o = n4246_o | n4248_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1249:33  */
  assign n4251_o = n3872_o == 12'b101100011100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1249:33  */
  assign n4252_o = n4249_o | n4251_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1249:56  */
  assign n4254_o = n3872_o == 12'b101100011101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1249:56  */
  assign n4255_o = n4252_o | n4254_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1249:79  */
  assign n4257_o = n3872_o == 12'b101100011110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1249:79  */
  assign n4258_o = n4255_o | n4257_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1249:102  */
  assign n4260_o = n3872_o == 12'b101100011111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1249:102  */
  assign n4261_o = n4258_o | n4260_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1249:125  */
  assign n4263_o = n3872_o == 12'b101110000011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1249:125  */
  assign n4264_o = n4261_o | n4263_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1250:33  */
  assign n4266_o = n3872_o == 12'b101110000100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1250:33  */
  assign n4267_o = n4264_o | n4266_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1250:56  */
  assign n4269_o = n3872_o == 12'b101110000101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1250:56  */
  assign n4270_o = n4267_o | n4269_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1250:79  */
  assign n4272_o = n3872_o == 12'b101110000110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1250:79  */
  assign n4273_o = n4270_o | n4272_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1250:102  */
  assign n4275_o = n3872_o == 12'b101110000111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1250:102  */
  assign n4276_o = n4273_o | n4275_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1250:125  */
  assign n4278_o = n3872_o == 12'b101110001000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1250:125  */
  assign n4279_o = n4276_o | n4278_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1250:148  */
  assign n4281_o = n3872_o == 12'b101110001001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1250:148  */
  assign n4282_o = n4279_o | n4281_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1251:33  */
  assign n4284_o = n3872_o == 12'b101110001010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1251:33  */
  assign n4285_o = n4282_o | n4284_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1251:56  */
  assign n4287_o = n3872_o == 12'b101110001011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1251:56  */
  assign n4288_o = n4285_o | n4287_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1251:79  */
  assign n4290_o = n3872_o == 12'b101110001100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1251:79  */
  assign n4291_o = n4288_o | n4290_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1251:102  */
  assign n4293_o = n3872_o == 12'b101110001101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1251:102  */
  assign n4294_o = n4291_o | n4293_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1251:125  */
  assign n4296_o = n3872_o == 12'b101110001110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1251:125  */
  assign n4297_o = n4294_o | n4296_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1251:148  */
  assign n4299_o = n3872_o == 12'b101110001111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1251:148  */
  assign n4300_o = n4297_o | n4299_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1252:33  */
  assign n4302_o = n3872_o == 12'b101110010000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1252:33  */
  assign n4303_o = n4300_o | n4302_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1252:56  */
  assign n4305_o = n3872_o == 12'b101110010001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1252:56  */
  assign n4306_o = n4303_o | n4305_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1252:79  */
  assign n4308_o = n3872_o == 12'b101110010010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1252:79  */
  assign n4309_o = n4306_o | n4308_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1252:102  */
  assign n4311_o = n3872_o == 12'b101110010011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1252:102  */
  assign n4312_o = n4309_o | n4311_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1252:125  */
  assign n4314_o = n3872_o == 12'b101110010100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1252:125  */
  assign n4315_o = n4312_o | n4314_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1252:148  */
  assign n4317_o = n3872_o == 12'b101110010101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1252:148  */
  assign n4318_o = n4315_o | n4317_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1253:33  */
  assign n4320_o = n3872_o == 12'b101110010110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1253:33  */
  assign n4321_o = n4318_o | n4320_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1253:56  */
  assign n4323_o = n3872_o == 12'b101110010111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1253:56  */
  assign n4324_o = n4321_o | n4323_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1253:79  */
  assign n4326_o = n3872_o == 12'b101110011000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1253:79  */
  assign n4327_o = n4324_o | n4326_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1253:102  */
  assign n4329_o = n3872_o == 12'b101110011001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1253:102  */
  assign n4330_o = n4327_o | n4329_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1253:125  */
  assign n4332_o = n3872_o == 12'b101110011010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1253:125  */
  assign n4333_o = n4330_o | n4332_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1253:148  */
  assign n4335_o = n3872_o == 12'b101110011011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1253:148  */
  assign n4336_o = n4333_o | n4335_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1254:33  */
  assign n4338_o = n3872_o == 12'b101110011100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1254:33  */
  assign n4339_o = n4336_o | n4338_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1254:56  */
  assign n4341_o = n3872_o == 12'b101110011101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1254:56  */
  assign n4342_o = n4339_o | n4341_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1254:79  */
  assign n4344_o = n3872_o == 12'b101110011110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1254:79  */
  assign n4345_o = n4342_o | n4344_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1254:102  */
  assign n4347_o = n3872_o == 12'b101110011111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1254:102  */
  assign n4348_o = n4345_o | n4347_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1254:125  */
  assign n4350_o = n3872_o == 12'b001100100011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1254:125  */
  assign n4351_o = n4348_o | n4350_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1255:33  */
  assign n4353_o = n3872_o == 12'b001100100100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1255:33  */
  assign n4354_o = n4351_o | n4353_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1255:56  */
  assign n4356_o = n3872_o == 12'b001100100101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1255:56  */
  assign n4357_o = n4354_o | n4356_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1255:79  */
  assign n4359_o = n3872_o == 12'b001100100110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1255:79  */
  assign n4360_o = n4357_o | n4359_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1255:102  */
  assign n4362_o = n3872_o == 12'b001100100111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1255:102  */
  assign n4363_o = n4360_o | n4362_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1255:125  */
  assign n4365_o = n3872_o == 12'b001100101000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1255:125  */
  assign n4366_o = n4363_o | n4365_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1255:148  */
  assign n4368_o = n3872_o == 12'b001100101001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1255:148  */
  assign n4369_o = n4366_o | n4368_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1256:33  */
  assign n4371_o = n3872_o == 12'b001100101010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1256:33  */
  assign n4372_o = n4369_o | n4371_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1256:56  */
  assign n4374_o = n3872_o == 12'b001100101011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1256:56  */
  assign n4375_o = n4372_o | n4374_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1256:79  */
  assign n4377_o = n3872_o == 12'b001100101100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1256:79  */
  assign n4378_o = n4375_o | n4377_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1256:102  */
  assign n4380_o = n3872_o == 12'b001100101101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1256:102  */
  assign n4381_o = n4378_o | n4380_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1256:125  */
  assign n4383_o = n3872_o == 12'b001100101110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1256:125  */
  assign n4384_o = n4381_o | n4383_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1256:148  */
  assign n4386_o = n3872_o == 12'b001100101111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1256:148  */
  assign n4387_o = n4384_o | n4386_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1257:33  */
  assign n4389_o = n3872_o == 12'b001100110000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1257:33  */
  assign n4390_o = n4387_o | n4389_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1257:56  */
  assign n4392_o = n3872_o == 12'b001100110001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1257:56  */
  assign n4393_o = n4390_o | n4392_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1257:79  */
  assign n4395_o = n3872_o == 12'b001100110010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1257:79  */
  assign n4396_o = n4393_o | n4395_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1257:102  */
  assign n4398_o = n3872_o == 12'b001100110011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1257:102  */
  assign n4399_o = n4396_o | n4398_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1257:125  */
  assign n4401_o = n3872_o == 12'b001100110100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1257:125  */
  assign n4402_o = n4399_o | n4401_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1257:148  */
  assign n4404_o = n3872_o == 12'b001100110101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1257:148  */
  assign n4405_o = n4402_o | n4404_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1258:33  */
  assign n4407_o = n3872_o == 12'b001100110110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1258:33  */
  assign n4408_o = n4405_o | n4407_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1258:56  */
  assign n4410_o = n3872_o == 12'b001100110111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1258:56  */
  assign n4411_o = n4408_o | n4410_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1258:79  */
  assign n4413_o = n3872_o == 12'b001100111000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1258:79  */
  assign n4414_o = n4411_o | n4413_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1258:102  */
  assign n4416_o = n3872_o == 12'b001100111001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1258:102  */
  assign n4417_o = n4414_o | n4416_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1258:125  */
  assign n4419_o = n3872_o == 12'b001100111010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1258:125  */
  assign n4420_o = n4417_o | n4419_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1258:148  */
  assign n4422_o = n3872_o == 12'b001100111011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1258:148  */
  assign n4423_o = n4420_o | n4422_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1259:33  */
  assign n4425_o = n3872_o == 12'b001100111100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1259:33  */
  assign n4426_o = n4423_o | n4425_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1259:56  */
  assign n4428_o = n3872_o == 12'b001100111101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1259:56  */
  assign n4429_o = n4426_o | n4428_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1259:79  */
  assign n4431_o = n3872_o == 12'b001100111110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1259:79  */
  assign n4432_o = n4429_o | n4431_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1259:102  */
  assign n4434_o = n3872_o == 12'b001100111111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1259:102  */
  assign n4435_o = n4432_o | n4434_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1263:7  */
  assign n4438_o = n3872_o == 12'b110000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1263:25  */
  assign n4440_o = n3872_o == 12'b101100000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1263:25  */
  assign n4441_o = n4438_o | n4440_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1263:41  */
  assign n4443_o = n3872_o == 12'b110000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1263:41  */
  assign n4444_o = n4441_o | n4443_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1263:55  */
  assign n4446_o = n3872_o == 12'b110000000010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1263:55  */
  assign n4447_o = n4444_o | n4446_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1263:72  */
  assign n4449_o = n3872_o == 12'b101100000010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1263:72  */
  assign n4450_o = n4447_o | n4449_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1263:90  */
  assign n4452_o = n3872_o == 12'b110010000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1263:90  */
  assign n4453_o = n4450_o | n4452_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1264:25  */
  assign n4455_o = n3872_o == 12'b101110000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1264:25  */
  assign n4456_o = n4453_o | n4455_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1264:41  */
  assign n4458_o = n3872_o == 12'b110010000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1264:41  */
  assign n4459_o = n4456_o | n4458_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1264:55  */
  assign n4461_o = n3872_o == 12'b110010000010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1264:55  */
  assign n4462_o = n4459_o | n4461_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1264:72  */
  assign n4464_o = n3872_o == 12'b101110000010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1264:72  */
  assign n4465_o = n4462_o | n4464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1268:7  */
  assign n4468_o = n3872_o == 12'b011110110000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1268:23  */
  assign n4470_o = n3872_o == 12'b011110110001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1268:23  */
  assign n4471_o = n4468_o | n4470_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1268:35  */
  assign n4473_o = n3872_o == 12'b011110110010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1268:35  */
  assign n4474_o = n4471_o | n4473_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1272:7  */
  assign n4477_o = n3872_o == 12'b011110100000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1272:26  */
  assign n4479_o = n3872_o == 12'b011110100001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1272:26  */
  assign n4480_o = n4477_o | n4479_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1272:41  */
  assign n4482_o = n3872_o == 12'b011110100010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1272:41  */
  assign n4483_o = n4480_o | n4482_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1272:56  */
  assign n4485_o = n3872_o == 12'b011110100011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1272:56  */
  assign n4486_o = n4483_o | n4485_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1272:71  */
  assign n4488_o = n3872_o == 12'b011110100100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1272:71  */
  assign n4489_o = n4486_o | n4488_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1272:85  */
  assign n4491_o = n3872_o == 12'b011110100101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1272:85  */
  assign n4492_o = n4489_o | n4491_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1272:102  */
  assign n4494_o = n3872_o == 12'b011110101000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1272:102  */
  assign n4495_o = n4492_o | n4494_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1272:119  */
  assign n4497_o = n3872_o == 12'b011110101010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1272:119  */
  assign n4498_o = n4495_o | n4497_o;
  assign n4499_o = {n4498_o, n4474_o, n4465_o, n4435_o, n4000_o, n3940_o, n3881_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1216:5  */
  always @*
    case (n4499_o)
      7'b1000000: n4508_o = 1'b0;
      7'b0100000: n4508_o = 1'b0;
      7'b0010000: n4508_o = 1'b1;
      7'b0001000: n4508_o = 1'b0;
      7'b0000100: n4508_o = 1'b0;
      7'b0000010: n4508_o = 1'b1;
      7'b0000001: n4508_o = 1'b0;
      default: n4508_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1287:17  */
  assign n4512_o = csr[11:10];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1287:32  */
  assign n4514_o = n4512_o == 2'b11;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1289:30  */
  assign n4515_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1289:77  */
  assign n4517_o = n4515_o == 3'b001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1290:30  */
  assign n4518_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1290:77  */
  assign n4520_o = n4518_o == 3'b101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1289:95  */
  assign n4521_o = n4517_o | n4520_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1291:21  */
  assign n4522_o = decode_aux[6];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1291:30  */
  assign n4523_o = ~n4522_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1290:96  */
  assign n4524_o = n4521_o | n4523_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1287:40  */
  assign n4525_o = n4514_o & n4524_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1287:5  */
  assign n4528_o = n4525_o ? 1'b0 : 1'b1;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1311:20  */
  assign n4547_o = csr[9:8];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1311:33  */
  assign n4549_o = n4547_o != 2'b00;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1311:51  */
  assign n4550_o = csr[121];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1311:65  */
  assign n4551_o = ~n4550_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1311:42  */
  assign n4552_o = n4549_o & n4551_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1311:5  */
  assign n4555_o = n4552_o ? 1'b0 : 1'b1;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1327:30  */
  assign n4558_o = execute_engine[22:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1329:7  */
  assign n4560_o = n4558_o == 7'b0110111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1329:25  */
  assign n4562_o = n4558_o == 7'b0010111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1329:25  */
  assign n4563_o = n4560_o | n4562_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1329:42  */
  assign n4565_o = n4558_o == 7'b1101111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1329:42  */
  assign n4566_o = n4563_o | n4565_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1335:34  */
  assign n4567_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1336:11  */
  assign n4569_o = n4567_o == 3'b000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1335:9  */
  always @*
    case (n4569_o)
      1'b1: n4572_o = 1'b0;
      default: n4572_o = 1'b1;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1333:7  */
  assign n4574_o = n4558_o == 7'b1100111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1342:34  */
  assign n4575_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1343:11  */
  assign n4577_o = n4575_o == 3'b000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1343:29  */
  assign n4579_o = n4575_o == 3'b001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1343:29  */
  assign n4580_o = n4577_o | n4579_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1343:44  */
  assign n4582_o = n4575_o == 3'b100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1343:44  */
  assign n4583_o = n4580_o | n4582_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1343:59  */
  assign n4585_o = n4575_o == 3'b101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1343:59  */
  assign n4586_o = n4583_o | n4585_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1343:74  */
  assign n4588_o = n4575_o == 3'b110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1343:74  */
  assign n4589_o = n4586_o | n4588_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1343:90  */
  assign n4591_o = n4575_o == 3'b111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1343:90  */
  assign n4592_o = n4589_o | n4591_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1342:9  */
  always @*
    case (n4592_o)
      1'b1: n4595_o = 1'b0;
      default: n4595_o = 1'b1;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1340:7  */
  assign n4597_o = n4558_o == 7'b1100011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1349:34  */
  assign n4598_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1350:11  */
  assign n4600_o = n4598_o == 3'b000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1350:28  */
  assign n4602_o = n4598_o == 3'b001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1350:28  */
  assign n4603_o = n4600_o | n4602_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1350:42  */
  assign n4605_o = n4598_o == 3'b010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1350:42  */
  assign n4606_o = n4603_o | n4605_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1350:56  */
  assign n4608_o = n4598_o == 3'b100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1350:56  */
  assign n4609_o = n4606_o | n4608_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1350:71  */
  assign n4611_o = n4598_o == 3'b101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1350:71  */
  assign n4612_o = n4609_o | n4611_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1349:9  */
  always @*
    case (n4612_o)
      1'b1: n4615_o = 1'b0;
      default: n4615_o = 1'b1;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1347:7  */
  assign n4617_o = n4558_o == 7'b0000011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1356:34  */
  assign n4618_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1357:11  */
  assign n4620_o = n4618_o == 3'b000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1357:28  */
  assign n4622_o = n4618_o == 3'b001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1357:28  */
  assign n4623_o = n4620_o | n4622_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1357:42  */
  assign n4625_o = n4618_o == 3'b010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1357:42  */
  assign n4626_o = n4623_o | n4625_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1356:9  */
  always @*
    case (n4626_o)
      1'b1: n4629_o = 1'b0;
      default: n4629_o = 1'b1;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1354:7  */
  assign n4631_o = n4558_o == 7'b0100011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1363:36  */
  assign n4632_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1363:83  */
  assign n4634_o = n4632_o == 3'b000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1363:126  */
  assign n4635_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1363:173  */
  assign n4637_o = n4635_o == 3'b101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1363:102  */
  assign n4638_o = n4634_o | n4637_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1364:35  */
  assign n4639_o = execute_engine[45:41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1364:84  */
  assign n4641_o = n4639_o == 5'b00000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1363:189  */
  assign n4642_o = n4638_o & n4641_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1364:120  */
  assign n4643_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1364:141  */
  assign n4644_o = ~n4643_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1364:95  */
  assign n4645_o = n4642_o & n4644_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1365:36  */
  assign n4646_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1365:83  */
  assign n4648_o = n4646_o == 3'b001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1366:36  */
  assign n4649_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1366:83  */
  assign n4651_o = n4649_o == 3'b010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1365:99  */
  assign n4652_o = n4648_o | n4651_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1367:36  */
  assign n4653_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1367:83  */
  assign n4655_o = n4653_o == 3'b011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1366:99  */
  assign n4656_o = n4652_o | n4655_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1368:36  */
  assign n4657_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1368:83  */
  assign n4659_o = n4657_o == 3'b100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1367:100  */
  assign n4660_o = n4656_o | n4659_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1369:36  */
  assign n4661_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1369:83  */
  assign n4663_o = n4661_o == 3'b110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1368:99  */
  assign n4664_o = n4660_o | n4663_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1370:36  */
  assign n4665_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1370:83  */
  assign n4667_o = n4665_o == 3'b111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1369:98  */
  assign n4668_o = n4664_o | n4667_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1371:36  */
  assign n4669_o = execute_engine[47:41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1371:83  */
  assign n4671_o = n4669_o == 7'b0000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1370:100  */
  assign n4672_o = n4668_o & n4671_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1364:149  */
  assign n4673_o = n4645_o | n4672_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1372:100  */
  assign n4674_o = decode_aux[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1372:84  */
  assign n4676_o = 1'b1 & n4674_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1371:98  */
  assign n4677_o = n4673_o | n4676_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1373:60  */
  assign n4678_o = decode_aux[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1373:44  */
  assign n4680_o = 1'b1 & n4678_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1372:117  */
  assign n4681_o = n4677_o | n4680_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1373:77  */
  assign n4683_o = n4681_o | 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1374:77  */
  assign n4685_o = n4683_o | 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1363:9  */
  assign n4688_o = n4685_o ? 1'b0 : 1'b1;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1361:7  */
  assign n4690_o = n4558_o == 7'b0110011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1383:34  */
  assign n4691_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1383:81  */
  assign n4693_o = n4691_o == 3'b000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1384:34  */
  assign n4694_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1384:81  */
  assign n4696_o = n4694_o == 3'b010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1383:100  */
  assign n4697_o = n4693_o | n4696_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1385:34  */
  assign n4698_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1385:81  */
  assign n4700_o = n4698_o == 3'b011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1384:97  */
  assign n4701_o = n4697_o | n4700_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1386:34  */
  assign n4702_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1386:81  */
  assign n4704_o = n4702_o == 3'b100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1385:98  */
  assign n4705_o = n4701_o | n4704_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1387:34  */
  assign n4706_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1387:81  */
  assign n4708_o = n4706_o == 3'b110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1386:97  */
  assign n4709_o = n4705_o | n4708_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1388:34  */
  assign n4710_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1388:81  */
  assign n4712_o = n4710_o == 3'b111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1387:96  */
  assign n4713_o = n4709_o | n4712_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1389:35  */
  assign n4714_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1389:82  */
  assign n4716_o = n4714_o == 3'b001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1390:35  */
  assign n4717_o = execute_engine[47:41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1390:82  */
  assign n4719_o = n4717_o == 7'b0000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1389:98  */
  assign n4720_o = n4716_o & n4719_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1388:97  */
  assign n4721_o = n4713_o | n4720_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1391:35  */
  assign n4722_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1391:82  */
  assign n4724_o = n4722_o == 3'b101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1392:36  */
  assign n4725_o = execute_engine[45:41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1392:85  */
  assign n4727_o = n4725_o == 5'b00000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1392:121  */
  assign n4728_o = execute_engine[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1392:142  */
  assign n4729_o = ~n4728_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1392:96  */
  assign n4730_o = n4727_o & n4729_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1391:97  */
  assign n4731_o = n4724_o & n4730_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1390:96  */
  assign n4732_o = n4721_o | n4731_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1392:152  */
  assign n4734_o = n4732_o | 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1383:9  */
  assign n4737_o = n4734_o ? 1'b0 : 1'b1;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1381:7  */
  assign n4739_o = n4558_o == 7'b0010011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1401:34  */
  assign n4740_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1402:11  */
  assign n4742_o = n4740_o == 3'b000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1403:11  */
  assign n4745_o = n4740_o == 3'b001;
  assign n4746_o = {n4745_o, n4742_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1401:9  */
  always @*
    case (n4746_o)
      2'b10: n4750_o = 1'b1;
      2'b01: n4750_o = 1'b0;
      default: n4750_o = 1'b1;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1399:7  */
  assign n4752_o = n4558_o == 7'b0001111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1409:33  */
  assign n4753_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1409:80  */
  assign n4755_o = n4753_o == 3'b000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1410:26  */
  assign n4756_o = decode_aux[6];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1410:58  */
  assign n4757_o = decode_aux[7];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1410:42  */
  assign n4758_o = n4756_o & n4757_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1411:38  */
  assign n4759_o = execute_engine[47:36];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1412:15  */
  assign n4761_o = n4759_o == 12'b000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1412:36  */
  assign n4763_o = n4759_o == 12'b000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1412:36  */
  assign n4764_o = n4761_o | n4763_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1413:81  */
  assign n4765_o = csr[120];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1413:73  */
  assign n4766_o = ~n4765_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1413:15  */
  assign n4768_o = n4759_o == 12'b001100000010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1414:82  */
  assign n4769_o = csr[120];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1414:74  */
  assign n4770_o = ~n4769_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1414:101  */
  assign n4771_o = csr[84];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1414:93  */
  assign n4772_o = n4770_o & n4771_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1414:15  */
  assign n4774_o = n4759_o == 12'b000100000101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1415:88  */
  assign n4775_o = debug_ctrl[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1415:73  */
  assign n4776_o = ~n4775_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1415:15  */
  assign n4778_o = n4759_o == 12'b011110110010;
  assign n4779_o = {n4778_o, n4774_o, n4768_o, n4764_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1411:13  */
  always @*
    case (n4779_o)
      4'b1000: n4782_o = n4776_o;
      4'b0100: n4782_o = n4772_o;
      4'b0010: n4782_o = n4766_o;
      4'b0001: n4782_o = 1'b0;
      default: n4782_o = 1'b1;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1410:11  */
  assign n4784_o = n4758_o ? n4782_o : 1'b1;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1421:30  */
  assign n4785_o = ~csr_reg_valid;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1421:54  */
  assign n4786_o = ~csr_rw_valid;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1421:37  */
  assign n4787_o = n4785_o | n4786_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1421:80  */
  assign n4788_o = ~csr_priv_valid;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1421:61  */
  assign n4789_o = n4787_o | n4788_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1422:36  */
  assign n4790_o = execute_engine[30:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1422:83  */
  assign n4792_o = n4790_o == 3'b100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1421:87  */
  assign n4793_o = n4789_o | n4792_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1421:9  */
  assign n4796_o = n4793_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1409:9  */
  assign n4797_o = n4755_o ? n4784_o : n4796_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1407:7  */
  assign n4799_o = n4558_o == 7'b1110011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1430:93  */
  assign n4801_o = decode_aux[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1430:78  */
  assign n4802_o = ~n4801_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1430:74  */
  assign n4804_o = 1'b1 | n4802_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1428:7  */
  assign n4806_o = n4558_o == 7'b1010011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1432:7  */
  assign n4809_o = n4558_o == 7'b0001011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1432:27  */
  assign n4811_o = n4558_o == 7'b0101011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1432:27  */
  assign n4812_o = n4809_o | n4811_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1432:44  */
  assign n4814_o = n4558_o == 7'b1011011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1432:44  */
  assign n4815_o = n4812_o | n4814_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1432:61  */
  assign n4817_o = n4558_o == 7'b1111011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1432:61  */
  assign n4818_o = n4815_o | n4817_o;
  assign n4819_o = {n4818_o, n4806_o, n4799_o, n4752_o, n4739_o, n4690_o, n4631_o, n4617_o, n4597_o, n4574_o, n4566_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1327:5  */
  always @*
    case (n4819_o)
      11'b10000000000: n4823_o = 1'b1;
      11'b01000000000: n4823_o = n4804_o;
      11'b00100000000: n4823_o = n4797_o;
      11'b00010000000: n4823_o = n4750_o;
      11'b00001000000: n4823_o = n4737_o;
      11'b00000100000: n4823_o = n4688_o;
      11'b00000010000: n4823_o = n4629_o;
      11'b00000001000: n4823_o = n4615_o;
      11'b00000000100: n4823_o = n4595_o;
      11'b00000000010: n4823_o = n4572_o;
      11'b00000000001: n4823_o = 1'b0;
      default: n4823_o = 1'b1;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1447:37  */
  assign n4826_o = illegal_cmd | alu_exc_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1448:85  */
  assign n4828_o = execute_engine[82];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1448:66  */
  assign n4830_o = 1'b1 & n4828_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1447:50  */
  assign n4831_o = n4826_o | n4830_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1449:47  */
  assign n4832_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1449:53  */
  assign n4834_o = n4832_o == 4'b0101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1449:83  */
  assign n4835_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1449:89  */
  assign n4837_o = n4835_o == 4'b0110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1449:64  */
  assign n4838_o = n4834_o | n4837_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1449:25  */
  assign n4839_o = n4838_o ? n4831_o : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1460:16  */
  assign n4842_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1473:60  */
  assign n4847_o = trap_ctrl[6];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1473:75  */
  assign n4848_o = n4847_o | ma_load_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1473:117  */
  assign n4849_o = trap_ctrl[95];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1473:103  */
  assign n4850_o = ~n4849_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1473:98  */
  assign n4851_o = n4848_o & n4850_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1474:60  */
  assign n4852_o = trap_ctrl[5];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1474:75  */
  assign n4853_o = n4852_o | ma_store_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1474:117  */
  assign n4854_o = trap_ctrl[95];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1474:103  */
  assign n4855_o = ~n4854_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1474:98  */
  assign n4856_o = n4853_o & n4855_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1475:60  */
  assign n4857_o = trap_ctrl[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1475:88  */
  assign n4858_o = trap_ctrl[98];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1475:75  */
  assign n4859_o = n4857_o | n4858_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1475:117  */
  assign n4860_o = trap_ctrl[95];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1475:103  */
  assign n4861_o = ~n4860_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1475:98  */
  assign n4862_o = n4859_o & n4861_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1478:61  */
  assign n4863_o = trap_ctrl[8];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1478:77  */
  assign n4864_o = n4863_o | be_load_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1478:119  */
  assign n4865_o = trap_ctrl[95];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1478:105  */
  assign n4866_o = ~n4865_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1478:100  */
  assign n4867_o = n4864_o & n4866_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1479:61  */
  assign n4868_o = trap_ctrl[7];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1479:77  */
  assign n4869_o = n4868_o | be_store_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1479:119  */
  assign n4870_o = trap_ctrl[95];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1479:105  */
  assign n4871_o = ~n4870_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1479:100  */
  assign n4872_o = n4869_o & n4871_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1480:61  */
  assign n4873_o = trap_ctrl[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1480:90  */
  assign n4874_o = trap_ctrl[97];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1480:77  */
  assign n4875_o = n4873_o | n4874_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1480:119  */
  assign n4876_o = trap_ctrl[95];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1480:105  */
  assign n4877_o = ~n4876_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1480:100  */
  assign n4878_o = n4875_o & n4877_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1483:62  */
  assign n4879_o = trap_ctrl[3];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1483:92  */
  assign n4880_o = trap_ctrl[100];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1483:79  */
  assign n4881_o = n4879_o | n4880_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1483:121  */
  assign n4882_o = trap_ctrl[95];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1483:107  */
  assign n4883_o = ~n4882_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1483:102  */
  assign n4884_o = n4881_o & n4883_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1484:62  */
  assign n4885_o = trap_ctrl[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1484:92  */
  assign n4886_o = trap_ctrl[99];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1484:79  */
  assign n4887_o = n4885_o | n4886_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1484:121  */
  assign n4888_o = trap_ctrl[95];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1484:107  */
  assign n4889_o = ~n4888_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1484:102  */
  assign n4890_o = n4887_o & n4889_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1493:61  */
  assign n4891_o = trap_ctrl[4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1493:88  */
  assign n4892_o = trap_ctrl[101];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1493:75  */
  assign n4893_o = n4891_o | n4892_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1493:100  */
  assign n4894_o = n4893_o | hw_trigger_fire;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1493:139  */
  assign n4895_o = trap_ctrl[95];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1493:125  */
  assign n4896_o = ~n4895_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1493:120  */
  assign n4897_o = n4894_o & n4896_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:64  */
  assign n4900_o = trap_ctrl[15];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:102  */
  assign n4901_o = csr[104];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:81  */
  assign n4902_o = n4900_o & n4901_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:116  */
  assign n4903_o = firq_i[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:107  */
  assign n4904_o = n4902_o | n4903_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:64  */
  assign n4905_o = trap_ctrl[16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:102  */
  assign n4906_o = csr[105];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:81  */
  assign n4907_o = n4905_o & n4906_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:116  */
  assign n4908_o = firq_i[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:107  */
  assign n4909_o = n4907_o | n4908_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:64  */
  assign n4910_o = trap_ctrl[17];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:102  */
  assign n4911_o = csr[106];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:81  */
  assign n4912_o = n4910_o & n4911_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:116  */
  assign n4913_o = firq_i[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:107  */
  assign n4914_o = n4912_o | n4913_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:64  */
  assign n4915_o = trap_ctrl[18];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:102  */
  assign n4916_o = csr[107];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:81  */
  assign n4917_o = n4915_o & n4916_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:116  */
  assign n4918_o = firq_i[3];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:107  */
  assign n4919_o = n4917_o | n4918_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:64  */
  assign n4920_o = trap_ctrl[19];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:102  */
  assign n4921_o = csr[108];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:81  */
  assign n4922_o = n4920_o & n4921_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:116  */
  assign n4923_o = firq_i[4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:107  */
  assign n4924_o = n4922_o | n4923_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:64  */
  assign n4925_o = trap_ctrl[20];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:102  */
  assign n4926_o = csr[109];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:81  */
  assign n4927_o = n4925_o & n4926_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:116  */
  assign n4928_o = firq_i[5];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:107  */
  assign n4929_o = n4927_o | n4928_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:64  */
  assign n4930_o = trap_ctrl[21];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:102  */
  assign n4931_o = csr[110];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:81  */
  assign n4932_o = n4930_o & n4931_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:116  */
  assign n4933_o = firq_i[6];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:107  */
  assign n4934_o = n4932_o | n4933_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:64  */
  assign n4935_o = trap_ctrl[22];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:102  */
  assign n4936_o = csr[111];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:81  */
  assign n4937_o = n4935_o & n4936_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:116  */
  assign n4938_o = firq_i[7];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:107  */
  assign n4939_o = n4937_o | n4938_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:64  */
  assign n4940_o = trap_ctrl[23];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:102  */
  assign n4941_o = csr[112];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:81  */
  assign n4942_o = n4940_o & n4941_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:116  */
  assign n4943_o = firq_i[8];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:107  */
  assign n4944_o = n4942_o | n4943_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:64  */
  assign n4945_o = trap_ctrl[24];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:102  */
  assign n4946_o = csr[113];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:81  */
  assign n4947_o = n4945_o & n4946_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:116  */
  assign n4948_o = firq_i[9];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:107  */
  assign n4949_o = n4947_o | n4948_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:64  */
  assign n4950_o = trap_ctrl[25];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:102  */
  assign n4951_o = csr[114];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:81  */
  assign n4952_o = n4950_o & n4951_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:116  */
  assign n4953_o = firq_i[10];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:107  */
  assign n4954_o = n4952_o | n4953_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:64  */
  assign n4955_o = trap_ctrl[26];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:102  */
  assign n4956_o = csr[115];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:81  */
  assign n4957_o = n4955_o & n4956_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:116  */
  assign n4958_o = firq_i[11];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:107  */
  assign n4959_o = n4957_o | n4958_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:64  */
  assign n4960_o = trap_ctrl[27];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:102  */
  assign n4961_o = csr[116];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:81  */
  assign n4962_o = n4960_o & n4961_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:116  */
  assign n4963_o = firq_i[12];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:107  */
  assign n4964_o = n4962_o | n4963_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:64  */
  assign n4965_o = trap_ctrl[28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:102  */
  assign n4966_o = csr[117];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:81  */
  assign n4967_o = n4965_o & n4966_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:116  */
  assign n4968_o = firq_i[13];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:107  */
  assign n4969_o = n4967_o | n4968_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:64  */
  assign n4970_o = trap_ctrl[29];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:102  */
  assign n4971_o = csr[118];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:81  */
  assign n4972_o = n4970_o & n4971_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:116  */
  assign n4973_o = firq_i[14];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:107  */
  assign n4974_o = n4972_o | n4973_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:64  */
  assign n4975_o = trap_ctrl[30];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:102  */
  assign n4976_o = csr[119];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:81  */
  assign n4977_o = n4975_o & n4976_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:116  */
  assign n4978_o = firq_i[15];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1518:107  */
  assign n4979_o = n4977_o | n4978_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1533:61  */
  assign n4982_o = trap_ctrl[12];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1533:85  */
  assign n4983_o = csr[85];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1533:77  */
  assign n4984_o = n4982_o & n4983_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1533:108  */
  assign n4985_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1533:139  */
  assign n4986_o = trap_ctrl[33];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1533:118  */
  assign n4987_o = n4985_o & n4986_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1533:94  */
  assign n4988_o = n4984_o | n4987_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1534:61  */
  assign n4989_o = trap_ctrl[14];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1534:85  */
  assign n4990_o = csr[86];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1534:77  */
  assign n4991_o = n4989_o & n4990_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1534:108  */
  assign n4992_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1534:139  */
  assign n4993_o = trap_ctrl[35];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1534:118  */
  assign n4994_o = n4992_o & n4993_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1534:94  */
  assign n4995_o = n4991_o | n4994_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1535:61  */
  assign n4996_o = trap_ctrl[13];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1535:85  */
  assign n4997_o = csr[87];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1535:77  */
  assign n4998_o = n4996_o & n4997_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1535:108  */
  assign n4999_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1535:139  */
  assign n5000_o = trap_ctrl[34];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1535:118  */
  assign n5001_o = n4999_o & n5000_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1535:94  */
  assign n5002_o = n4998_o | n5001_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:64  */
  assign n5003_o = trap_ctrl[15];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:97  */
  assign n5004_o = csr[88];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:81  */
  assign n5005_o = n5003_o & n5004_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:116  */
  assign n5006_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:147  */
  assign n5007_o = trap_ctrl[36];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:126  */
  assign n5008_o = n5006_o & n5007_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:102  */
  assign n5009_o = n5005_o | n5008_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:64  */
  assign n5010_o = trap_ctrl[16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:97  */
  assign n5011_o = csr[89];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:81  */
  assign n5012_o = n5010_o & n5011_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:116  */
  assign n5013_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:147  */
  assign n5014_o = trap_ctrl[37];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:126  */
  assign n5015_o = n5013_o & n5014_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:102  */
  assign n5016_o = n5012_o | n5015_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:64  */
  assign n5017_o = trap_ctrl[17];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:97  */
  assign n5018_o = csr[90];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:81  */
  assign n5019_o = n5017_o & n5018_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:116  */
  assign n5020_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:147  */
  assign n5021_o = trap_ctrl[38];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:126  */
  assign n5022_o = n5020_o & n5021_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:102  */
  assign n5023_o = n5019_o | n5022_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:64  */
  assign n5024_o = trap_ctrl[18];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:97  */
  assign n5025_o = csr[91];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:81  */
  assign n5026_o = n5024_o & n5025_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:116  */
  assign n5027_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:147  */
  assign n5028_o = trap_ctrl[39];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:126  */
  assign n5029_o = n5027_o & n5028_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:102  */
  assign n5030_o = n5026_o | n5029_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:64  */
  assign n5031_o = trap_ctrl[19];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:97  */
  assign n5032_o = csr[92];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:81  */
  assign n5033_o = n5031_o & n5032_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:116  */
  assign n5034_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:147  */
  assign n5035_o = trap_ctrl[40];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:126  */
  assign n5036_o = n5034_o & n5035_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:102  */
  assign n5037_o = n5033_o | n5036_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:64  */
  assign n5038_o = trap_ctrl[20];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:97  */
  assign n5039_o = csr[93];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:81  */
  assign n5040_o = n5038_o & n5039_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:116  */
  assign n5041_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:147  */
  assign n5042_o = trap_ctrl[41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:126  */
  assign n5043_o = n5041_o & n5042_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:102  */
  assign n5044_o = n5040_o | n5043_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:64  */
  assign n5045_o = trap_ctrl[21];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:97  */
  assign n5046_o = csr[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:81  */
  assign n5047_o = n5045_o & n5046_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:116  */
  assign n5048_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:147  */
  assign n5049_o = trap_ctrl[42];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:126  */
  assign n5050_o = n5048_o & n5049_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:102  */
  assign n5051_o = n5047_o | n5050_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:64  */
  assign n5052_o = trap_ctrl[22];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:97  */
  assign n5053_o = csr[95];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:81  */
  assign n5054_o = n5052_o & n5053_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:116  */
  assign n5055_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:147  */
  assign n5056_o = trap_ctrl[43];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:126  */
  assign n5057_o = n5055_o & n5056_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:102  */
  assign n5058_o = n5054_o | n5057_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:64  */
  assign n5059_o = trap_ctrl[23];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:97  */
  assign n5060_o = csr[96];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:81  */
  assign n5061_o = n5059_o & n5060_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:116  */
  assign n5062_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:147  */
  assign n5063_o = trap_ctrl[44];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:126  */
  assign n5064_o = n5062_o & n5063_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:102  */
  assign n5065_o = n5061_o | n5064_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:64  */
  assign n5066_o = trap_ctrl[24];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:97  */
  assign n5067_o = csr[97];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:81  */
  assign n5068_o = n5066_o & n5067_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:116  */
  assign n5069_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:147  */
  assign n5070_o = trap_ctrl[45];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:126  */
  assign n5071_o = n5069_o & n5070_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:102  */
  assign n5072_o = n5068_o | n5071_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:64  */
  assign n5073_o = trap_ctrl[25];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:97  */
  assign n5074_o = csr[98];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:81  */
  assign n5075_o = n5073_o & n5074_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:116  */
  assign n5076_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:147  */
  assign n5077_o = trap_ctrl[46];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:126  */
  assign n5078_o = n5076_o & n5077_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:102  */
  assign n5079_o = n5075_o | n5078_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:64  */
  assign n5080_o = trap_ctrl[26];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:97  */
  assign n5081_o = csr[99];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:81  */
  assign n5082_o = n5080_o & n5081_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:116  */
  assign n5083_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:147  */
  assign n5084_o = trap_ctrl[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:126  */
  assign n5085_o = n5083_o & n5084_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:102  */
  assign n5086_o = n5082_o | n5085_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:64  */
  assign n5087_o = trap_ctrl[27];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:97  */
  assign n5088_o = csr[100];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:81  */
  assign n5089_o = n5087_o & n5088_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:116  */
  assign n5090_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:147  */
  assign n5091_o = trap_ctrl[48];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:126  */
  assign n5092_o = n5090_o & n5091_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:102  */
  assign n5093_o = n5089_o | n5092_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:64  */
  assign n5094_o = trap_ctrl[28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:97  */
  assign n5095_o = csr[101];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:81  */
  assign n5096_o = n5094_o & n5095_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:116  */
  assign n5097_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:147  */
  assign n5098_o = trap_ctrl[49];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:126  */
  assign n5099_o = n5097_o & n5098_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:102  */
  assign n5100_o = n5096_o | n5099_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:64  */
  assign n5101_o = trap_ctrl[29];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:97  */
  assign n5102_o = csr[102];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:81  */
  assign n5103_o = n5101_o & n5102_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:116  */
  assign n5104_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:147  */
  assign n5105_o = trap_ctrl[50];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:126  */
  assign n5106_o = n5104_o & n5105_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:102  */
  assign n5107_o = n5103_o | n5106_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:64  */
  assign n5108_o = trap_ctrl[30];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:97  */
  assign n5109_o = csr[103];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:81  */
  assign n5110_o = n5108_o & n5109_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:116  */
  assign n5111_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:147  */
  assign n5112_o = trap_ctrl[51];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:126  */
  assign n5113_o = n5111_o & n5112_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1539:102  */
  assign n5114_o = n5110_o | n5113_o;
  assign n5117_o = {1'b0, 1'b0, n4867_o, n4872_o, n4851_o, n4856_o, n4897_o, n4884_o, n4862_o, n4890_o, n4878_o};
  assign n5118_o = {1'b0, 1'b0, n5114_o, n5107_o, n5100_o, n5093_o, n5086_o, n5079_o, n5072_o, n5065_o, n5058_o, n5051_o, n5044_o, n5037_o, n5030_o, n5023_o, n5016_o, n5009_o, n4995_o, n5002_o, n4988_o, 1'b0, 1'b0, n4979_o, n4974_o, n4969_o, n4964_o, n4959_o, n4954_o, n4949_o, n4944_o, n4939_o, n4934_o, n4929_o, n4924_o, n4919_o, n4914_o, n4909_o, n4904_o, mext_irq_i, mtime_irq_i, msw_irq_i};
  assign n5123_o = {21'b000000000000000000000, 21'b000000000000000000000};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1559:16  */
  assign n5128_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1562:21  */
  assign n5131_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1562:31  */
  assign n5132_o = ~n5131_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1563:24  */
  assign n5133_o = trap_ctrl[11];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1565:24  */
  assign n5134_o = trap_ctrl[54];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1565:61  */
  assign n5135_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1565:67  */
  assign n5137_o = n5135_o == 4'b0101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1565:97  */
  assign n5138_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1565:103  */
  assign n5140_o = n5138_o == 4'b0010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1565:78  */
  assign n5141_o = n5137_o | n5140_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1565:40  */
  assign n5142_o = n5134_o & n5141_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1563:41  */
  assign n5143_o = n5133_o | n5142_o;
  assign n5145_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1563:9  */
  assign n5146_o = n5143_o ? 1'b1 : n5145_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1569:23  */
  assign n5147_o = trap_ctrl[95];
  assign n5149_o = trap_ctrl[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1569:9  */
  assign n5150_o = n5147_o ? 1'b0 : n5149_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1562:7  */
  assign n5151_o = n5132_o ? n5146_o : n5150_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1580:57  */
  assign n5158_o = trap_ctrl[10:0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5164_o = n5158_o[10];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5166_o = 1'b0 | n5164_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5168_o = n5158_o[9];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5169_o = n5166_o | n5168_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5170_o = n5158_o[8];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5171_o = n5169_o | n5170_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5172_o = n5158_o[7];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5173_o = n5171_o | n5172_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5174_o = n5158_o[6];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5175_o = n5173_o | n5174_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5176_o = n5158_o[5];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5177_o = n5175_o | n5176_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5178_o = n5158_o[4];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5179_o = n5177_o | n5178_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5180_o = n5158_o[3];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5181_o = n5179_o | n5180_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5182_o = n5158_o[2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5183_o = n5181_o | n5182_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5184_o = n5158_o[1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5185_o = n5183_o | n5184_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5186_o = n5158_o[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5187_o = n5185_o | n5186_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1580:29  */
  assign n5188_o = n5187_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1585:36  */
  assign n5192_o = trap_ctrl[51:33];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5198_o = n5192_o[18];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5200_o = 1'b0 | n5198_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5202_o = n5192_o[17];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5203_o = n5200_o | n5202_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5204_o = n5192_o[16];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5205_o = n5203_o | n5204_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5206_o = n5192_o[15];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5207_o = n5205_o | n5206_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5208_o = n5192_o[14];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5209_o = n5207_o | n5208_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5210_o = n5192_o[13];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5211_o = n5209_o | n5210_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5212_o = n5192_o[12];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5213_o = n5211_o | n5212_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5214_o = n5192_o[11];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5215_o = n5213_o | n5214_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5216_o = n5192_o[10];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5217_o = n5215_o | n5216_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5218_o = n5192_o[9];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5219_o = n5217_o | n5218_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5220_o = n5192_o[8];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5221_o = n5219_o | n5220_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5222_o = n5192_o[7];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5223_o = n5221_o | n5222_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5224_o = n5192_o[6];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5225_o = n5223_o | n5224_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5226_o = n5192_o[5];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5227_o = n5225_o | n5226_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5228_o = n5192_o[4];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5229_o = n5227_o | n5228_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5230_o = n5192_o[3];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5231_o = n5229_o | n5230_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5232_o = n5192_o[2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5233_o = n5231_o | n5232_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5234_o = n5192_o[1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5235_o = n5233_o | n5234_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n5236_o = n5192_o[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n5237_o = n5235_o | n5236_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1586:12  */
  assign n5238_o = csr[80];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1586:39  */
  assign n5239_o = csr[120];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1586:49  */
  assign n5240_o = ~n5239_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1586:31  */
  assign n5241_o = n5238_o | n5240_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1585:81  */
  assign n5242_o = n5237_o & n5241_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1587:18  */
  assign n5243_o = debug_ctrl[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1587:26  */
  assign n5244_o = ~n5243_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1586:67  */
  assign n5245_o = n5242_o & n5244_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1588:11  */
  assign n5246_o = csr[330];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1588:21  */
  assign n5247_o = ~n5246_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1587:33  */
  assign n5248_o = n5245_o & n5247_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1590:23  */
  assign n5249_o = trap_ctrl[53];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1589:7  */
  assign n5250_o = n5248_o | n5249_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1591:23  */
  assign n5251_o = trap_ctrl[52];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1590:46  */
  assign n5252_o = n5250_o | n5251_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1583:29  */
  assign n5253_o = n5252_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1594:38  */
  assign n5255_o = execute_engine[116:86];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1594:56  */
  assign n5257_o = {n5255_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1594:86  */
  assign n5258_o = trap_ctrl[61];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1594:131  */
  assign n5259_o = trap_ctrl[61:55];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1594:137  */
  assign n5261_o = n5259_o == 7'b0000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1594:117  */
  assign n5262_o = n5258_o | n5261_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1594:63  */
  assign n5263_o = n5262_o ? n5257_o : n5266_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1595:43  */
  assign n5264_o = execute_engine[214:184];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1595:61  */
  assign n5266_o = {n5264_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1604:31  */
  assign n5269_o = trap_ctrl[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1605:31  */
  assign n5271_o = trap_ctrl[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1606:31  */
  assign n5273_o = trap_ctrl[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1607:31  */
  assign n5275_o = trap_ctrl[3];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1607:108  */
  assign n5276_o = csr[120];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1607:102  */
  assign n5278_o = {5'b00010, n5276_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1607:124  */
  assign n5279_o = csr[120];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1607:118  */
  assign n5280_o = {n5278_o, n5279_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1608:31  */
  assign n5281_o = trap_ctrl[4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1609:31  */
  assign n5283_o = trap_ctrl[5];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1610:31  */
  assign n5285_o = trap_ctrl[6];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1611:31  */
  assign n5287_o = trap_ctrl[7];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1612:31  */
  assign n5289_o = trap_ctrl[8];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1614:31  */
  assign n5291_o = trap_ctrl[52];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1615:31  */
  assign n5293_o = trap_ctrl[10];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1616:31  */
  assign n5295_o = trap_ctrl[9];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1617:31  */
  assign n5297_o = trap_ctrl[53];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1619:31  */
  assign n5299_o = trap_ctrl[36];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1620:31  */
  assign n5301_o = trap_ctrl[37];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1621:31  */
  assign n5303_o = trap_ctrl[38];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1622:31  */
  assign n5305_o = trap_ctrl[39];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1623:31  */
  assign n5307_o = trap_ctrl[40];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1624:31  */
  assign n5309_o = trap_ctrl[41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1625:31  */
  assign n5311_o = trap_ctrl[42];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1626:31  */
  assign n5313_o = trap_ctrl[43];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1627:31  */
  assign n5315_o = trap_ctrl[44];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1628:31  */
  assign n5317_o = trap_ctrl[45];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1629:31  */
  assign n5319_o = trap_ctrl[46];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1630:31  */
  assign n5321_o = trap_ctrl[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1631:31  */
  assign n5323_o = trap_ctrl[48];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1632:31  */
  assign n5325_o = trap_ctrl[49];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1633:31  */
  assign n5327_o = trap_ctrl[50];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1634:31  */
  assign n5329_o = trap_ctrl[51];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1636:31  */
  assign n5331_o = trap_ctrl[35];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1637:31  */
  assign n5333_o = trap_ctrl[33];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1637:7  */
  assign n5337_o = n5333_o ? 7'b1000011 : 7'b1000111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1636:7  */
  assign n5338_o = n5331_o ? 7'b1001011 : n5337_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1634:7  */
  assign n5339_o = n5329_o ? 7'b1011111 : n5338_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1633:7  */
  assign n5340_o = n5327_o ? 7'b1011110 : n5339_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1632:7  */
  assign n5341_o = n5325_o ? 7'b1011101 : n5340_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1631:7  */
  assign n5342_o = n5323_o ? 7'b1011100 : n5341_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1630:7  */
  assign n5343_o = n5321_o ? 7'b1011011 : n5342_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1629:7  */
  assign n5344_o = n5319_o ? 7'b1011010 : n5343_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1628:7  */
  assign n5345_o = n5317_o ? 7'b1011001 : n5344_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1627:7  */
  assign n5346_o = n5315_o ? 7'b1011000 : n5345_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1626:7  */
  assign n5347_o = n5313_o ? 7'b1010111 : n5346_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1625:7  */
  assign n5348_o = n5311_o ? 7'b1010110 : n5347_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1624:7  */
  assign n5349_o = n5309_o ? 7'b1010101 : n5348_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1623:7  */
  assign n5350_o = n5307_o ? 7'b1010100 : n5349_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1622:7  */
  assign n5351_o = n5305_o ? 7'b1010011 : n5350_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1621:7  */
  assign n5352_o = n5303_o ? 7'b1010010 : n5351_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1620:7  */
  assign n5353_o = n5301_o ? 7'b1010001 : n5352_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1619:7  */
  assign n5354_o = n5299_o ? 7'b1010000 : n5353_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1617:7  */
  assign n5355_o = n5297_o ? 7'b1100100 : n5354_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1616:7  */
  assign n5356_o = n5295_o ? 7'b0100001 : n5355_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1615:7  */
  assign n5357_o = n5293_o ? 7'b0100010 : n5356_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1614:7  */
  assign n5358_o = n5291_o ? 7'b1100011 : n5357_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1612:7  */
  assign n5359_o = n5289_o ? 7'b0000101 : n5358_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1611:7  */
  assign n5360_o = n5287_o ? 7'b0000111 : n5359_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1610:7  */
  assign n5361_o = n5285_o ? 7'b0000100 : n5360_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1609:7  */
  assign n5362_o = n5283_o ? 7'b0000110 : n5361_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1608:7  */
  assign n5363_o = n5281_o ? 7'b0000011 : n5362_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1607:7  */
  assign n5364_o = n5275_o ? n5280_o : n5363_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1606:7  */
  assign n5365_o = n5273_o ? 7'b0000010 : n5364_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1605:7  */
  assign n5366_o = n5271_o ? 7'b0000001 : n5365_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1604:7  */
  assign n5367_o = n5269_o ? 7'b0000000 : n5366_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1654:29  */
  assign n5373_o = execute_engine[30];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1656:48  */
  assign n5374_o = execute_engine[35:31];
  assign n5376_o = n5375_o[31:5];
  assign n5377_o = {n5376_o, n5374_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1654:5  */
  assign n5378_o = n5373_o ? n5377_o : rs1_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1661:30  */
  assign n5379_o = execute_engine[29:28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1662:39  */
  assign n5380_o = csr[79:48];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1662:45  */
  assign n5381_o = n5380_o | n5378_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1662:7  */
  assign n5383_o = n5379_o == 2'b10;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1663:39  */
  assign n5384_o = csr[79:48];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1663:50  */
  assign n5385_o = ~n5378_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1663:45  */
  assign n5386_o = n5384_o & n5385_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1663:7  */
  assign n5388_o = n5379_o == 2'b11;
  assign n5389_o = {n5388_o, n5383_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1661:5  */
  always @*
    case (n5389_o)
      2'b10: n5390_o = n5386_o;
      2'b01: n5390_o = n5381_o;
      default: n5390_o = n5378_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1673:16  */
  assign n5393_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1709:21  */
  assign n5427_o = csr[13];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1709:54  */
  assign n5428_o = trap_ctrl[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1709:33  */
  assign n5429_o = ~n5428_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1709:28  */
  assign n5430_o = n5427_o & n5429_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1717:15  */
  assign n5432_o = csr[12];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1736:21  */
  assign n5433_o = csr[11:3];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1736:35  */
  assign n5435_o = n5433_o == 9'b001100000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1738:23  */
  assign n5436_o = csr[2:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1738:36  */
  assign n5438_o = n5436_o == 3'b000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1739:42  */
  assign n5439_o = csr[19];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1740:42  */
  assign n5440_o = csr[23];
  assign n5441_o = {n5440_o, n5439_o};
  assign n5442_o = csr[81:80];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1736:9  */
  assign n5443_o = n5466_o ? n5441_o : n5442_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1748:23  */
  assign n5444_o = csr[2:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1748:36  */
  assign n5446_o = n5444_o == 3'b100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1749:38  */
  assign n5447_o = csr[19];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1750:38  */
  assign n5448_o = csr[23];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1751:38  */
  assign n5449_o = csr[27];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1752:38  */
  assign n5450_o = csr[47:32];
  assign n5451_o = {n5450_o, n5448_o, n5449_o, n5447_o};
  assign n5452_o = csr[103:85];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1736:9  */
  assign n5453_o = n5468_o ? n5451_o : n5452_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1755:23  */
  assign n5454_o = csr[2:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1755:36  */
  assign n5456_o = n5454_o == 3'b101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1756:35  */
  assign n5457_o = csr[47:18];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1756:53  */
  assign n5459_o = {n5457_o, 2'b00};
  assign n5460_o = csr[191:160];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1736:9  */
  assign n5461_o = n5470_o ? n5459_o : n5460_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1736:9  */
  assign n5466_o = n5435_o & n5438_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1736:9  */
  assign n5468_o = n5435_o & n5446_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1736:9  */
  assign n5470_o = n5435_o & n5456_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1774:21  */
  assign n5471_o = csr[11:4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1774:35  */
  assign n5473_o = n5471_o == 8'b00110100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1776:23  */
  assign n5474_o = csr[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1776:36  */
  assign n5476_o = n5474_o == 4'b0000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1777:33  */
  assign n5477_o = csr[47:16];
  assign n5478_o = csr[255:224];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1776:11  */
  assign n5479_o = n5476_o ? n5477_o : n5478_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1780:23  */
  assign n5480_o = csr[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1780:36  */
  assign n5482_o = n5480_o == 4'b0001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1781:29  */
  assign n5483_o = csr[47:16];
  assign n5484_o = csr[153:122];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1780:11  */
  assign n5485_o = n5482_o ? n5483_o : n5484_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1784:23  */
  assign n5486_o = csr[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1784:36  */
  assign n5488_o = n5486_o == 4'b0010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1785:36  */
  assign n5489_o = csr[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1785:52  */
  assign n5490_o = csr[20:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1785:41  */
  assign n5491_o = {n5489_o, n5490_o};
  assign n5492_o = csr[159:154];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1784:11  */
  assign n5493_o = n5488_o ? n5491_o : n5492_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1788:22  */
  assign n5494_o = csr[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1788:35  */
  assign n5496_o = n5494_o == 4'b0011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1789:29  */
  assign n5497_o = csr[47:16];
  assign n5498_o = csr[223:192];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1788:10  */
  assign n5499_o = n5496_o ? n5497_o : n5498_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1792:23  */
  assign n5500_o = csr[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1792:36  */
  assign n5502_o = n5500_o == 4'b0100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1793:43  */
  assign n5503_o = csr[47:32];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1774:9  */
  assign n5504_o = n5507_o ? n5503_o : 16'b1111111111111111;
  assign n5505_o = {n5493_o, n5485_o};
  assign n5506_o = {n5479_o, n5499_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1774:9  */
  assign n5507_o = n5473_o & n5502_o;
  assign n5508_o = csr[159:122];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1774:9  */
  assign n5509_o = n5473_o ? n5505_o : n5508_o;
  assign n5510_o = csr[255:192];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1774:9  */
  assign n5511_o = n5473_o ? n5506_o : n5510_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1799:21  */
  assign n5512_o = csr[11:5];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1799:35  */
  assign n5514_o = n5512_o == 7'b0011001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1801:23  */
  assign n5515_o = csr[4:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1801:36  */
  assign n5517_o = n5515_o == 5'b00000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1803:48  */
  assign n5518_o = csr[16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1804:48  */
  assign n5519_o = csr[18];
  assign n5520_o = csr[288];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1717:7  */
  assign n5521_o = n5601_o ? n5518_o : n5520_o;
  assign n5522_o = csr[290];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1717:7  */
  assign n5523_o = n5603_o ? n5519_o : n5522_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1799:9  */
  assign n5525_o = n5514_o & n5517_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1799:9  */
  assign n5527_o = n5514_o & n5517_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1871:23  */
  assign n5528_o = trap_ctrl[95];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1877:42  */
  assign n5529_o = trap_ctrl[61];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1877:82  */
  assign n5530_o = trap_ctrl[59:55];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1877:65  */
  assign n5531_o = {n5529_o, n5530_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1879:35  */
  assign n5532_o = trap_ctrl[93:62];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1881:28  */
  assign n5533_o = trap_ctrl[61:55];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1883:47  */
  assign n5534_o = execute_engine[116:86];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1883:65  */
  assign n5536_o = {n5534_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1882:15  */
  assign n5538_o = n5533_o == 7'b0000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1882:31  */
  assign n5540_o = n5533_o == 7'b0000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1882:31  */
  assign n5541_o = n5538_o | n5540_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1884:15  */
  assign n5543_o = n5533_o == 7'b0000100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1884:31  */
  assign n5545_o = n5533_o == 7'b0000101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1884:31  */
  assign n5546_o = n5543_o | n5545_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1884:44  */
  assign n5548_o = n5533_o == 7'b0000110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1884:44  */
  assign n5549_o = n5546_o | n5548_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1884:57  */
  assign n5551_o = n5533_o == 7'b0000111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1884:57  */
  assign n5552_o = n5549_o | n5551_o;
  assign n5554_o = {n5552_o, n5541_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1881:13  */
  always @*
    case (n5554_o)
      2'b10: n5555_o = mar_i;
      2'b01: n5555_o = n5536_o;
      default: n5555_o = 32'b00000000000000000000000000000000;
    endcase
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1892:37  */
  assign n5558_o = csr[80];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1893:37  */
  assign n5559_o = csr[120];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1910:26  */
  assign n5560_o = trap_ctrl[96];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1933:37  */
  assign n5563_o = csr[81];
  assign n5565_o = {1'b1, 1'b1, n5563_o};
  assign n5566_o = csr[82:80];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1910:9  */
  assign n5567_o = n5560_o ? n5565_o : n5566_o;
  assign n5568_o = csr[120];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1910:9  */
  assign n5569_o = n5560_o ? 1'b1 : n5568_o;
  assign n5570_o = {n5559_o, n5558_o, 1'b0};
  assign n5571_o = {n5531_o, n5532_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1871:9  */
  assign n5572_o = n5528_o ? n5570_o : n5567_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1871:9  */
  assign n5573_o = n5528_o ? 1'b1 : n5569_o;
  assign n5574_o = csr[159:122];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1871:9  */
  assign n5575_o = n5528_o ? n5571_o : n5574_o;
  assign n5576_o = csr[223:192];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1871:9  */
  assign n5577_o = n5528_o ? n5555_o : n5576_o;
  assign n5578_o = {n5504_o, n5453_o};
  assign n5579_o = {n5511_o, n5461_o, n5509_o};
  assign n5580_o = n5572_o[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1717:7  */
  assign n5581_o = n5432_o ? n5443_o : n5580_o;
  assign n5582_o = n5572_o[2];
  assign n5583_o = csr[82];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1717:7  */
  assign n5584_o = n5432_o ? n5583_o : n5582_o;
  assign n5585_o = csr[103:85];
  assign n5586_o = {16'b1111111111111111, n5585_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1717:7  */
  assign n5587_o = n5432_o ? n5578_o : n5586_o;
  assign n5588_o = csr[120];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1717:7  */
  assign n5589_o = n5432_o ? n5588_o : n5573_o;
  assign n5590_o = n5579_o[37:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1717:7  */
  assign n5591_o = n5432_o ? n5590_o : n5575_o;
  assign n5592_o = n5579_o[69:38];
  assign n5593_o = csr[191:160];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1717:7  */
  assign n5594_o = n5432_o ? n5592_o : n5593_o;
  assign n5595_o = n5579_o[101:70];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1717:7  */
  assign n5596_o = n5432_o ? n5595_o : n5577_o;
  assign n5597_o = n5579_o[133:102];
  assign n5598_o = csr[255:224];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1717:7  */
  assign n5599_o = n5432_o ? n5597_o : n5598_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1717:7  */
  assign n5601_o = n5432_o & n5525_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1717:7  */
  assign n5603_o = n5432_o & n5527_o;
  assign n5626_o = {n5589_o, n5587_o, 1'b0, 1'b0, n5584_o, n5581_o};
  assign n5627_o = {3'b000, 1'b1, 1'b0, 1'b0, 1'b0, 5'b00000, 3'b000, 29'b00000000000000000000000000000, n5523_o, 1'b0, n5521_o, 32'b00000000000000000000000000000000, n5599_o, n5596_o, n5594_o, n5591_o};
  assign n5628_o = {1'b0, 1'b0, 1'b0, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000};
  assign n5639_o = {1'b1, 16'b0000000000000000, 16'b0000000000000000, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
  assign n5640_o = {3'b000, 1'b1, 1'b0, 1'b0, 1'b0, 5'b00000, 3'b000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 32'b00011001100010000000011100000100, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 6'b000000, 32'b00000000000000000000000000000000};
  assign n5641_o = {1'b0, 1'b0, 1'b0, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2000:38  */
  assign n5650_o = 1'b0 ? 1'b1 : n5651_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2000:118  */
  assign n5651_o = csr[120];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2124:24  */
  assign n5705_o = csr[15];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2135:9  */
  assign n5708_o = csr_raddr == 12'b000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2138:9  */
  assign n5710_o = csr_raddr == 12'b000000000010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2141:9  */
  assign n5712_o = csr_raddr == 12'b000000000011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2147:32  */
  assign n5713_o = csr[80];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2148:32  */
  assign n5714_o = csr[81];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2149:53  */
  assign n5715_o = csr[82];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2149:53  */
  assign n5716_o = csr[82];
  assign n5717_o = {n5715_o, n5716_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2150:32  */
  assign n5718_o = csr[83];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2151:32  */
  assign n5719_o = csr[84];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2151:43  */
  assign n5722_o = n5719_o & 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2146:9  */
  assign n5724_o = csr_raddr == 12'b001100000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2156:9  */
  assign n5741_o = csr_raddr == 12'b001100000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2168:32  */
  assign n5742_o = csr[85];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2169:32  */
  assign n5743_o = csr[87];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2170:32  */
  assign n5744_o = csr[86];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2171:42  */
  assign n5745_o = csr[103:88];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2167:9  */
  assign n5747_o = csr_raddr == 12'b001100000100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2174:33  */
  assign n5748_o = csr[191:162];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2174:51  */
  assign n5750_o = {n5748_o, 2'b00};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2173:9  */
  assign n5752_o = csr_raddr == 12'b001100000101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2176:9  */
  assign n5754_o = csr_raddr == 12'b001100000110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2194:28  */
  assign n5755_o = csr[255:224];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2193:9  */
  assign n5757_o = csr_raddr == 12'b001101000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2197:32  */
  assign n5758_o = csr[153:123];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2197:50  */
  assign n5760_o = {n5758_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2196:9  */
  assign n5762_o = csr_raddr == 12'b001101000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2200:46  */
  assign n5763_o = csr[159];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2201:46  */
  assign n5764_o = csr[158:154];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2199:9  */
  assign n5766_o = csr_raddr == 12'b001101000010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2204:28  */
  assign n5767_o = csr[223:192];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2203:9  */
  assign n5769_o = csr_raddr == 12'b001101000011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2207:55  */
  assign n5770_o = trap_ctrl[12];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2208:55  */
  assign n5771_o = trap_ctrl[13];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2209:55  */
  assign n5772_o = trap_ctrl[14];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2210:55  */
  assign n5773_o = trap_ctrl[30:15];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2206:9  */
  assign n5775_o = csr_raddr == 12'b001101000100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2215:9  */
  assign n5777_o = csr_raddr == 12'b001110100000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2215:28  */
  assign n5779_o = csr_raddr == 12'b001110100001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2215:28  */
  assign n5780_o = n5777_o | n5779_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2215:44  */
  assign n5782_o = csr_raddr == 12'b001110100010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2215:44  */
  assign n5783_o = n5780_o | n5782_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2215:60  */
  assign n5785_o = csr_raddr == 12'b001110100011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2215:60  */
  assign n5786_o = n5783_o | n5785_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2219:9  */
  assign n5788_o = csr_raddr == 12'b001110110000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2219:30  */
  assign n5790_o = csr_raddr == 12'b001110110001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2219:30  */
  assign n5791_o = n5788_o | n5790_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2219:48  */
  assign n5793_o = csr_raddr == 12'b001110110010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2219:48  */
  assign n5794_o = n5791_o | n5793_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2219:66  */
  assign n5796_o = csr_raddr == 12'b001110110011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2219:66  */
  assign n5797_o = n5794_o | n5796_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2219:84  */
  assign n5799_o = csr_raddr == 12'b001110110100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2219:84  */
  assign n5800_o = n5797_o | n5799_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2220:30  */
  assign n5802_o = csr_raddr == 12'b001110110101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2220:30  */
  assign n5803_o = n5800_o | n5802_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2220:48  */
  assign n5805_o = csr_raddr == 12'b001110110110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2220:48  */
  assign n5806_o = n5803_o | n5805_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2220:66  */
  assign n5808_o = csr_raddr == 12'b001110110111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2220:66  */
  assign n5809_o = n5806_o | n5808_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2220:84  */
  assign n5811_o = csr_raddr == 12'b001110111000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2220:84  */
  assign n5812_o = n5809_o | n5811_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2221:30  */
  assign n5814_o = csr_raddr == 12'b001110111001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2221:30  */
  assign n5815_o = n5812_o | n5814_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2221:48  */
  assign n5817_o = csr_raddr == 12'b001110111010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2221:48  */
  assign n5818_o = n5815_o | n5817_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2221:66  */
  assign n5820_o = csr_raddr == 12'b001110111011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2221:66  */
  assign n5821_o = n5818_o | n5820_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2221:84  */
  assign n5823_o = csr_raddr == 12'b001110111100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2221:84  */
  assign n5824_o = n5821_o | n5823_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2222:30  */
  assign n5826_o = csr_raddr == 12'b001110111101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2222:30  */
  assign n5827_o = n5824_o | n5826_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2222:48  */
  assign n5829_o = csr_raddr == 12'b001110111110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2222:48  */
  assign n5830_o = n5827_o | n5829_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2222:66  */
  assign n5832_o = csr_raddr == 12'b001110111111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2222:66  */
  assign n5833_o = n5830_o | n5832_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2229:46  */
  assign n5834_o = csr[288];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2230:46  */
  assign n5835_o = csr[290];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2227:9  */
  assign n5837_o = csr_raddr == 12'b001100100000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2237:9  */
  assign n5839_o = csr_raddr == 12'b001100100011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2238:9  */
  assign n5841_o = csr_raddr == 12'b001100100100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2239:9  */
  assign n5843_o = csr_raddr == 12'b001100100101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2240:9  */
  assign n5845_o = csr_raddr == 12'b001100100110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2241:9  */
  assign n5847_o = csr_raddr == 12'b001100100111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2242:9  */
  assign n5849_o = csr_raddr == 12'b001100101000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2243:9  */
  assign n5851_o = csr_raddr == 12'b001100101001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2244:9  */
  assign n5853_o = csr_raddr == 12'b001100101010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2245:9  */
  assign n5855_o = csr_raddr == 12'b001100101011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2246:9  */
  assign n5857_o = csr_raddr == 12'b001100101100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2247:9  */
  assign n5859_o = csr_raddr == 12'b001100101101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2248:9  */
  assign n5861_o = csr_raddr == 12'b001100101110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2249:9  */
  assign n5863_o = csr_raddr == 12'b001100101111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2250:9  */
  assign n5865_o = csr_raddr == 12'b001100110000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2251:9  */
  assign n5867_o = csr_raddr == 12'b001100110001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2252:9  */
  assign n5869_o = csr_raddr == 12'b001100110010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2253:9  */
  assign n5871_o = csr_raddr == 12'b001100110011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2254:9  */
  assign n5873_o = csr_raddr == 12'b001100110100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2255:9  */
  assign n5875_o = csr_raddr == 12'b001100110101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2256:9  */
  assign n5877_o = csr_raddr == 12'b001100110110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2257:9  */
  assign n5879_o = csr_raddr == 12'b001100110111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2258:9  */
  assign n5881_o = csr_raddr == 12'b001100111000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2259:9  */
  assign n5883_o = csr_raddr == 12'b001100111001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2260:9  */
  assign n5885_o = csr_raddr == 12'b001100111010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2261:9  */
  assign n5887_o = csr_raddr == 12'b001100111011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2262:9  */
  assign n5889_o = csr_raddr == 12'b001100111100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2263:9  */
  assign n5891_o = csr_raddr == 12'b001100111101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2264:9  */
  assign n5893_o = csr_raddr == 12'b001100111110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2265:9  */
  assign n5895_o = csr_raddr == 12'b001100111111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2270:117  */
  assign n5896_o = cnt_lo_rd[1023:992];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2270:9  */
  assign n5898_o = csr_raddr == 12'b101100000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2270:34  */
  assign n5900_o = csr_raddr == 12'b110000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2270:34  */
  assign n5901_o = n5898_o | n5900_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2271:117  */
  assign n5902_o = cnt_lo_rd[991:960];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2271:9  */
  assign n5904_o = csr_raddr == 12'b101100000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2271:34  */
  assign n5906_o = csr_raddr == 12'b110000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2271:34  */
  assign n5907_o = n5904_o | n5906_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2272:117  */
  assign n5908_o = cnt_lo_rd[959:928];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2272:9  */
  assign n5910_o = csr_raddr == 12'b101100000010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2272:34  */
  assign n5912_o = csr_raddr == 12'b110000000010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2272:34  */
  assign n5913_o = n5910_o | n5912_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2273:9  */
  assign n5915_o = csr_raddr == 12'b101100000011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2273:34  */
  assign n5917_o = csr_raddr == 12'b110000000011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2273:34  */
  assign n5918_o = n5915_o | n5917_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2274:9  */
  assign n5920_o = csr_raddr == 12'b101100000100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2274:34  */
  assign n5922_o = csr_raddr == 12'b110000000100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2274:34  */
  assign n5923_o = n5920_o | n5922_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2275:9  */
  assign n5925_o = csr_raddr == 12'b101100000101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2275:34  */
  assign n5927_o = csr_raddr == 12'b110000000101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2275:34  */
  assign n5928_o = n5925_o | n5927_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2276:9  */
  assign n5930_o = csr_raddr == 12'b101100000110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2276:34  */
  assign n5932_o = csr_raddr == 12'b110000000110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2276:34  */
  assign n5933_o = n5930_o | n5932_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2277:9  */
  assign n5935_o = csr_raddr == 12'b101100000111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2277:34  */
  assign n5937_o = csr_raddr == 12'b110000000111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2277:34  */
  assign n5938_o = n5935_o | n5937_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2278:9  */
  assign n5940_o = csr_raddr == 12'b101100001000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2278:34  */
  assign n5942_o = csr_raddr == 12'b110000001000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2278:34  */
  assign n5943_o = n5940_o | n5942_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2279:9  */
  assign n5945_o = csr_raddr == 12'b101100001001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2279:34  */
  assign n5947_o = csr_raddr == 12'b110000001001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2279:34  */
  assign n5948_o = n5945_o | n5947_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2280:9  */
  assign n5950_o = csr_raddr == 12'b101100001010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2280:34  */
  assign n5952_o = csr_raddr == 12'b110000001010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2280:34  */
  assign n5953_o = n5950_o | n5952_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2281:9  */
  assign n5955_o = csr_raddr == 12'b101100001011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2281:34  */
  assign n5957_o = csr_raddr == 12'b110000001011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2281:34  */
  assign n5958_o = n5955_o | n5957_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2282:9  */
  assign n5960_o = csr_raddr == 12'b101100001100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2282:34  */
  assign n5962_o = csr_raddr == 12'b110000001100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2282:34  */
  assign n5963_o = n5960_o | n5962_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2283:9  */
  assign n5965_o = csr_raddr == 12'b101100001101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2283:34  */
  assign n5967_o = csr_raddr == 12'b110000001101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2283:34  */
  assign n5968_o = n5965_o | n5967_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2284:9  */
  assign n5970_o = csr_raddr == 12'b101100001110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2284:34  */
  assign n5972_o = csr_raddr == 12'b110000001110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2284:34  */
  assign n5973_o = n5970_o | n5972_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2285:9  */
  assign n5975_o = csr_raddr == 12'b101100001111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2285:34  */
  assign n5977_o = csr_raddr == 12'b110000001111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2285:34  */
  assign n5978_o = n5975_o | n5977_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2286:9  */
  assign n5980_o = csr_raddr == 12'b101100010000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2286:34  */
  assign n5982_o = csr_raddr == 12'b110000010000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2286:34  */
  assign n5983_o = n5980_o | n5982_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2287:9  */
  assign n5985_o = csr_raddr == 12'b101100010001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2287:34  */
  assign n5987_o = csr_raddr == 12'b110000010001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2287:34  */
  assign n5988_o = n5985_o | n5987_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2288:9  */
  assign n5990_o = csr_raddr == 12'b101100010010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2288:34  */
  assign n5992_o = csr_raddr == 12'b110000010010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2288:34  */
  assign n5993_o = n5990_o | n5992_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2289:9  */
  assign n5995_o = csr_raddr == 12'b101100010011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2289:34  */
  assign n5997_o = csr_raddr == 12'b110000010011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2289:34  */
  assign n5998_o = n5995_o | n5997_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2290:9  */
  assign n6000_o = csr_raddr == 12'b101100010100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2290:34  */
  assign n6002_o = csr_raddr == 12'b110000010100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2290:34  */
  assign n6003_o = n6000_o | n6002_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2291:9  */
  assign n6005_o = csr_raddr == 12'b101100010101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2291:34  */
  assign n6007_o = csr_raddr == 12'b110000010101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2291:34  */
  assign n6008_o = n6005_o | n6007_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2292:9  */
  assign n6010_o = csr_raddr == 12'b101100010110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2292:34  */
  assign n6012_o = csr_raddr == 12'b110000010110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2292:34  */
  assign n6013_o = n6010_o | n6012_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2293:9  */
  assign n6015_o = csr_raddr == 12'b101100010111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2293:34  */
  assign n6017_o = csr_raddr == 12'b110000010111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2293:34  */
  assign n6018_o = n6015_o | n6017_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2294:9  */
  assign n6020_o = csr_raddr == 12'b101100011000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2294:34  */
  assign n6022_o = csr_raddr == 12'b110000011000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2294:34  */
  assign n6023_o = n6020_o | n6022_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2295:9  */
  assign n6025_o = csr_raddr == 12'b101100011001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2295:34  */
  assign n6027_o = csr_raddr == 12'b110000011001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2295:34  */
  assign n6028_o = n6025_o | n6027_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2296:9  */
  assign n6030_o = csr_raddr == 12'b101100011010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2296:34  */
  assign n6032_o = csr_raddr == 12'b110000011010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2296:34  */
  assign n6033_o = n6030_o | n6032_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2297:9  */
  assign n6035_o = csr_raddr == 12'b101100011011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2297:34  */
  assign n6037_o = csr_raddr == 12'b110000011011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2297:34  */
  assign n6038_o = n6035_o | n6037_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2298:9  */
  assign n6040_o = csr_raddr == 12'b101100011100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2298:34  */
  assign n6042_o = csr_raddr == 12'b110000011100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2298:34  */
  assign n6043_o = n6040_o | n6042_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2299:9  */
  assign n6045_o = csr_raddr == 12'b101100011101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2299:34  */
  assign n6047_o = csr_raddr == 12'b110000011101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2299:34  */
  assign n6048_o = n6045_o | n6047_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2300:9  */
  assign n6050_o = csr_raddr == 12'b101100011110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2300:34  */
  assign n6052_o = csr_raddr == 12'b110000011110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2300:34  */
  assign n6053_o = n6050_o | n6052_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2301:9  */
  assign n6055_o = csr_raddr == 12'b101100011111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2301:34  */
  assign n6057_o = csr_raddr == 12'b110000011111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2301:34  */
  assign n6058_o = n6055_o | n6057_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2304:119  */
  assign n6059_o = cnt_hi_rd[1023:992];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2304:9  */
  assign n6061_o = csr_raddr == 12'b101110000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2304:35  */
  assign n6063_o = csr_raddr == 12'b110010000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2304:35  */
  assign n6064_o = n6061_o | n6063_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2305:119  */
  assign n6065_o = cnt_hi_rd[991:960];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2305:9  */
  assign n6067_o = csr_raddr == 12'b101110000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2305:35  */
  assign n6069_o = csr_raddr == 12'b110010000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2305:35  */
  assign n6070_o = n6067_o | n6069_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2306:119  */
  assign n6071_o = cnt_hi_rd[959:928];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2306:9  */
  assign n6073_o = csr_raddr == 12'b101110000010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2306:35  */
  assign n6075_o = csr_raddr == 12'b110010000010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2306:35  */
  assign n6076_o = n6073_o | n6075_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2307:9  */
  assign n6078_o = csr_raddr == 12'b101110000011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2307:35  */
  assign n6080_o = csr_raddr == 12'b110010000011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2307:35  */
  assign n6081_o = n6078_o | n6080_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2308:9  */
  assign n6083_o = csr_raddr == 12'b101110000100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2308:35  */
  assign n6085_o = csr_raddr == 12'b110010000100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2308:35  */
  assign n6086_o = n6083_o | n6085_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2309:9  */
  assign n6088_o = csr_raddr == 12'b101110000101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2309:35  */
  assign n6090_o = csr_raddr == 12'b110010000101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2309:35  */
  assign n6091_o = n6088_o | n6090_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2310:9  */
  assign n6093_o = csr_raddr == 12'b101110000110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2310:35  */
  assign n6095_o = csr_raddr == 12'b110010000110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2310:35  */
  assign n6096_o = n6093_o | n6095_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2311:9  */
  assign n6098_o = csr_raddr == 12'b101110000111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2311:35  */
  assign n6100_o = csr_raddr == 12'b110010000111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2311:35  */
  assign n6101_o = n6098_o | n6100_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2312:9  */
  assign n6103_o = csr_raddr == 12'b101110001000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2312:35  */
  assign n6105_o = csr_raddr == 12'b110010001000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2312:35  */
  assign n6106_o = n6103_o | n6105_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2313:9  */
  assign n6108_o = csr_raddr == 12'b101110001001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2313:35  */
  assign n6110_o = csr_raddr == 12'b110010001001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2313:35  */
  assign n6111_o = n6108_o | n6110_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2314:9  */
  assign n6113_o = csr_raddr == 12'b101110001010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2314:35  */
  assign n6115_o = csr_raddr == 12'b110010001010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2314:35  */
  assign n6116_o = n6113_o | n6115_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2315:9  */
  assign n6118_o = csr_raddr == 12'b101110001011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2315:35  */
  assign n6120_o = csr_raddr == 12'b110010001011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2315:35  */
  assign n6121_o = n6118_o | n6120_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2316:9  */
  assign n6123_o = csr_raddr == 12'b101110001100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2316:35  */
  assign n6125_o = csr_raddr == 12'b110010001100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2316:35  */
  assign n6126_o = n6123_o | n6125_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2317:9  */
  assign n6128_o = csr_raddr == 12'b101110001101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2317:35  */
  assign n6130_o = csr_raddr == 12'b110010001101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2317:35  */
  assign n6131_o = n6128_o | n6130_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2318:9  */
  assign n6133_o = csr_raddr == 12'b101110001110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2318:35  */
  assign n6135_o = csr_raddr == 12'b110010001110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2318:35  */
  assign n6136_o = n6133_o | n6135_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2319:9  */
  assign n6138_o = csr_raddr == 12'b101110001111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2319:35  */
  assign n6140_o = csr_raddr == 12'b110010001111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2319:35  */
  assign n6141_o = n6138_o | n6140_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2320:9  */
  assign n6143_o = csr_raddr == 12'b101110010000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2320:35  */
  assign n6145_o = csr_raddr == 12'b110010010000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2320:35  */
  assign n6146_o = n6143_o | n6145_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2321:9  */
  assign n6148_o = csr_raddr == 12'b101110010001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2321:35  */
  assign n6150_o = csr_raddr == 12'b110010010001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2321:35  */
  assign n6151_o = n6148_o | n6150_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2322:9  */
  assign n6153_o = csr_raddr == 12'b101110010010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2322:35  */
  assign n6155_o = csr_raddr == 12'b110010010010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2322:35  */
  assign n6156_o = n6153_o | n6155_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2323:9  */
  assign n6158_o = csr_raddr == 12'b101110010011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2323:35  */
  assign n6160_o = csr_raddr == 12'b110010010011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2323:35  */
  assign n6161_o = n6158_o | n6160_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2324:9  */
  assign n6163_o = csr_raddr == 12'b101110010100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2324:35  */
  assign n6165_o = csr_raddr == 12'b110010010100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2324:35  */
  assign n6166_o = n6163_o | n6165_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2325:9  */
  assign n6168_o = csr_raddr == 12'b101110010101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2325:35  */
  assign n6170_o = csr_raddr == 12'b110010010101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2325:35  */
  assign n6171_o = n6168_o | n6170_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2326:9  */
  assign n6173_o = csr_raddr == 12'b101110010110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2326:35  */
  assign n6175_o = csr_raddr == 12'b110010010110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2326:35  */
  assign n6176_o = n6173_o | n6175_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2327:9  */
  assign n6178_o = csr_raddr == 12'b101110010111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2327:35  */
  assign n6180_o = csr_raddr == 12'b110010010111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2327:35  */
  assign n6181_o = n6178_o | n6180_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2328:9  */
  assign n6183_o = csr_raddr == 12'b101110011000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2328:35  */
  assign n6185_o = csr_raddr == 12'b110010011000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2328:35  */
  assign n6186_o = n6183_o | n6185_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2329:9  */
  assign n6188_o = csr_raddr == 12'b101110011001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2329:35  */
  assign n6190_o = csr_raddr == 12'b110010011001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2329:35  */
  assign n6191_o = n6188_o | n6190_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2330:9  */
  assign n6193_o = csr_raddr == 12'b101110011010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2330:35  */
  assign n6195_o = csr_raddr == 12'b110010011010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2330:35  */
  assign n6196_o = n6193_o | n6195_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2331:9  */
  assign n6198_o = csr_raddr == 12'b101110011011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2331:35  */
  assign n6200_o = csr_raddr == 12'b110010011011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2331:35  */
  assign n6201_o = n6198_o | n6200_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2332:9  */
  assign n6203_o = csr_raddr == 12'b101110011100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2332:35  */
  assign n6205_o = csr_raddr == 12'b110010011100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2332:35  */
  assign n6206_o = n6203_o | n6205_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2333:9  */
  assign n6208_o = csr_raddr == 12'b101110011101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2333:35  */
  assign n6210_o = csr_raddr == 12'b110010011101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2333:35  */
  assign n6211_o = n6208_o | n6210_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2334:9  */
  assign n6213_o = csr_raddr == 12'b101110011110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2334:35  */
  assign n6215_o = csr_raddr == 12'b110010011110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2334:35  */
  assign n6216_o = n6213_o | n6215_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2335:9  */
  assign n6218_o = csr_raddr == 12'b101110011111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2335:35  */
  assign n6220_o = csr_raddr == 12'b110010011111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2335:35  */
  assign n6221_o = n6218_o | n6220_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2339:9  */
  assign n6224_o = csr_raddr == 12'b111100010001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2340:9  */
  assign n6227_o = csr_raddr == 12'b111100010010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2341:9  */
  assign n6230_o = csr_raddr == 12'b111100010011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2342:9  */
  assign n6233_o = csr_raddr == 12'b111100010100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2347:9  */
  assign n6235_o = csr_raddr == 12'b011110110000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2348:9  */
  assign n6237_o = csr_raddr == 12'b011110110001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2349:9  */
  assign n6239_o = csr_raddr == 12'b011110110010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2354:9  */
  assign n6241_o = csr_raddr == 12'b011110100001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2355:9  */
  assign n6243_o = csr_raddr == 12'b011110100010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2357:9  */
  assign n6245_o = csr_raddr == 12'b011110100100;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2365:9  */
  assign n6274_o = csr_raddr == 12'b111111000000;
  assign n6276_o = {n6274_o, n6245_o, n6243_o, n6241_o, n6239_o, n6237_o, n6235_o, n6233_o, n6230_o, n6227_o, n6224_o, n6221_o, n6216_o, n6211_o, n6206_o, n6201_o, n6196_o, n6191_o, n6186_o, n6181_o, n6176_o, n6171_o, n6166_o, n6161_o, n6156_o, n6151_o, n6146_o, n6141_o, n6136_o, n6131_o, n6126_o, n6121_o, n6116_o, n6111_o, n6106_o, n6101_o, n6096_o, n6091_o, n6086_o, n6081_o, n6076_o, n6070_o, n6064_o, n6058_o, n6053_o, n6048_o, n6043_o, n6038_o, n6033_o, n6028_o, n6023_o, n6018_o, n6013_o, n6008_o, n6003_o, n5998_o, n5993_o, n5988_o, n5983_o, n5978_o, n5973_o, n5968_o, n5963_o, n5958_o, n5953_o, n5948_o, n5943_o, n5938_o, n5933_o, n5928_o, n5923_o, n5918_o, n5913_o, n5907_o, n5901_o, n5895_o, n5893_o, n5891_o, n5889_o, n5887_o, n5885_o, n5883_o, n5881_o, n5879_o, n5877_o, n5875_o, n5873_o, n5871_o, n5869_o, n5867_o, n5865_o, n5863_o, n5861_o, n5859_o, n5857_o, n5855_o, n5853_o, n5851_o, n5849_o, n5847_o, n5845_o, n5843_o, n5841_o, n5839_o, n5837_o, n5833_o, n5786_o, n5775_o, n5769_o, n5766_o, n5762_o, n5757_o, n5754_o, n5752_o, n5747_o, n5741_o, n5724_o, n5712_o, n5710_o, n5708_o};
  assign n6277_o = n5750_o[0];
  assign n6278_o = n5755_o[0];
  assign n6279_o = n5760_o[0];
  assign n6280_o = n5764_o[0];
  assign n6281_o = n5767_o[0];
  assign n6282_o = n5896_o[0];
  assign n6283_o = n5902_o[0];
  assign n6284_o = n5908_o[0];
  assign n6285_o = n6059_o[0];
  assign n6286_o = n6065_o[0];
  assign n6287_o = n6071_o[0];
  assign n6288_o = n6222_o[0];
  assign n6289_o = n6225_o[0];
  assign n6290_o = n6228_o[0];
  assign n6291_o = n6231_o[0];
  assign n6292_o = n6275_o[0];
  assign n6293_o = n5706_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = 1'b1;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6291_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6290_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6289_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6288_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6287_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6286_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6285_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6294_o = n6284_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6294_o = n6283_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6294_o = n6282_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6294_o = n5834_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6294_o = n6281_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6294_o = n6280_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6294_o = n6279_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6294_o = n6278_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6294_o = n6277_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6294_o = n6293_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6294_o = n6293_o;
      default: n6294_o = n6292_o;
    endcase
  assign n6295_o = n5750_o[1];
  assign n6296_o = n5755_o[1];
  assign n6297_o = n5760_o[1];
  assign n6298_o = n5764_o[1];
  assign n6299_o = n5767_o[1];
  assign n6300_o = n5896_o[1];
  assign n6301_o = n5902_o[1];
  assign n6302_o = n5908_o[1];
  assign n6303_o = n6059_o[1];
  assign n6304_o = n6065_o[1];
  assign n6305_o = n6071_o[1];
  assign n6306_o = n6222_o[1];
  assign n6307_o = n6225_o[1];
  assign n6308_o = n6228_o[1];
  assign n6309_o = n6231_o[1];
  assign n6310_o = n6275_o[1];
  assign n6311_o = n5706_o[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = 1'b0;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6309_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6308_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6307_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6306_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6305_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6304_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6303_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6312_o = n6302_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6312_o = n6301_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6312_o = n6300_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6312_o = n6299_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6312_o = n6298_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6312_o = n6297_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6312_o = n6296_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6312_o = n6295_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6312_o = 1'b0;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6312_o = n6311_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6312_o = n6311_o;
      default: n6312_o = n6310_o;
    endcase
  assign n6313_o = n5750_o[2];
  assign n6314_o = n5755_o[2];
  assign n6315_o = n5760_o[2];
  assign n6316_o = n5764_o[2];
  assign n6317_o = n5767_o[2];
  assign n6318_o = n5896_o[2];
  assign n6319_o = n5902_o[2];
  assign n6320_o = n5908_o[2];
  assign n6321_o = n6059_o[2];
  assign n6322_o = n6065_o[2];
  assign n6323_o = n6071_o[2];
  assign n6324_o = n6222_o[2];
  assign n6325_o = n6225_o[2];
  assign n6326_o = n6228_o[2];
  assign n6327_o = n6231_o[2];
  assign n6328_o = n6275_o[2];
  assign n6329_o = n5706_o[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = 1'b0;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6327_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6326_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6325_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6324_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6323_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6322_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6321_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6330_o = n6320_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6330_o = n6319_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6330_o = n6318_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6330_o = n5835_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6330_o = n6317_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6330_o = n6316_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6330_o = n6315_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6330_o = n6314_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6330_o = n6313_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6330_o = 1'b1;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6330_o = n6329_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6330_o = n6329_o;
      default: n6330_o = n6328_o;
    endcase
  assign n6331_o = n5750_o[3];
  assign n6332_o = n5755_o[3];
  assign n6333_o = n5760_o[3];
  assign n6334_o = n5764_o[3];
  assign n6335_o = n5767_o[3];
  assign n6336_o = n5896_o[3];
  assign n6337_o = n5902_o[3];
  assign n6338_o = n5908_o[3];
  assign n6339_o = n6059_o[3];
  assign n6340_o = n6065_o[3];
  assign n6341_o = n6071_o[3];
  assign n6342_o = n6222_o[3];
  assign n6343_o = n6225_o[3];
  assign n6344_o = n6228_o[3];
  assign n6345_o = n6231_o[3];
  assign n6346_o = n6275_o[3];
  assign n6347_o = n5706_o[3];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = 1'b0;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6345_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6344_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6343_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6342_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6341_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6340_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6339_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6348_o = n6338_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6348_o = n6337_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6348_o = n6336_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6348_o = n5770_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6348_o = n6335_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6348_o = n6334_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6348_o = n6333_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6348_o = n6332_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6348_o = n6331_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6348_o = n5742_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6348_o = n5713_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6348_o = n6347_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6348_o = n6347_o;
      default: n6348_o = n6346_o;
    endcase
  assign n6349_o = n5750_o[4];
  assign n6350_o = n5755_o[4];
  assign n6351_o = n5760_o[4];
  assign n6352_o = n5764_o[4];
  assign n6353_o = n5767_o[4];
  assign n6354_o = n5896_o[4];
  assign n6355_o = n5902_o[4];
  assign n6356_o = n5908_o[4];
  assign n6357_o = n6059_o[4];
  assign n6358_o = n6065_o[4];
  assign n6359_o = n6071_o[4];
  assign n6360_o = n6222_o[4];
  assign n6361_o = n6225_o[4];
  assign n6362_o = n6228_o[4];
  assign n6363_o = n6231_o[4];
  assign n6364_o = n6275_o[4];
  assign n6365_o = n5706_o[4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = 1'b0;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6363_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6362_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6361_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6360_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6359_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6358_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6357_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6366_o = n6356_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6366_o = n6355_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6366_o = n6354_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6366_o = n6353_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6366_o = n6352_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6366_o = n6351_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6366_o = n6350_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6366_o = n6349_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6366_o = 1'b0;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6366_o = n6365_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6366_o = n6365_o;
      default: n6366_o = n6364_o;
    endcase
  assign n6367_o = n5750_o[5];
  assign n6368_o = n5755_o[5];
  assign n6369_o = n5760_o[5];
  assign n6370_o = n5767_o[5];
  assign n6371_o = n5896_o[5];
  assign n6372_o = n5902_o[5];
  assign n6373_o = n5908_o[5];
  assign n6374_o = n6059_o[5];
  assign n6375_o = n6065_o[5];
  assign n6376_o = n6071_o[5];
  assign n6377_o = n6222_o[5];
  assign n6378_o = n6228_o[5];
  assign n6379_o = n6231_o[5];
  assign n6380_o = n6275_o[5];
  assign n6381_o = n5706_o[5];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = 1'b0;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6379_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6378_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6377_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6376_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6375_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6374_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6382_o = n6373_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6382_o = n6372_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6382_o = n6371_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6382_o = n6370_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6382_o = n6369_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6382_o = n6368_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6382_o = n6367_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6382_o = n6381_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6382_o = n6381_o;
      default: n6382_o = n6380_o;
    endcase
  assign n6383_o = n5750_o[6];
  assign n6384_o = n5755_o[6];
  assign n6385_o = n5760_o[6];
  assign n6386_o = n5767_o[6];
  assign n6387_o = n5896_o[6];
  assign n6388_o = n5902_o[6];
  assign n6389_o = n5908_o[6];
  assign n6390_o = n6059_o[6];
  assign n6391_o = n6065_o[6];
  assign n6392_o = n6071_o[6];
  assign n6393_o = n6222_o[6];
  assign n6394_o = n6228_o[6];
  assign n6395_o = n6231_o[6];
  assign n6396_o = n6275_o[6];
  assign n6397_o = n5706_o[6];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6395_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6394_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6393_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6392_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6391_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6390_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6398_o = n6389_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6398_o = n6388_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6398_o = n6387_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6398_o = n6386_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6398_o = n6385_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6398_o = n6384_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6398_o = n6383_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6398_o = n6397_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6398_o = n6397_o;
      default: n6398_o = n6396_o;
    endcase
  assign n6399_o = n5750_o[7];
  assign n6400_o = n5755_o[7];
  assign n6401_o = n5760_o[7];
  assign n6402_o = n5767_o[7];
  assign n6403_o = n5896_o[7];
  assign n6404_o = n5902_o[7];
  assign n6405_o = n5908_o[7];
  assign n6406_o = n6059_o[7];
  assign n6407_o = n6065_o[7];
  assign n6408_o = n6071_o[7];
  assign n6409_o = n6222_o[7];
  assign n6410_o = n6228_o[7];
  assign n6411_o = n6231_o[7];
  assign n6412_o = n6275_o[7];
  assign n6413_o = n5706_o[7];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = 1'b1;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6411_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6410_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6409_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6408_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6407_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6406_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6414_o = n6405_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6414_o = n6404_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6414_o = n6403_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6414_o = n5771_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6414_o = n6402_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6414_o = n6401_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6414_o = n6400_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6414_o = n6399_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6414_o = n5743_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6414_o = n5714_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6414_o = n6413_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6414_o = n6413_o;
      default: n6414_o = n6412_o;
    endcase
  assign n6415_o = n5750_o[8];
  assign n6416_o = n5755_o[8];
  assign n6417_o = n5760_o[8];
  assign n6418_o = n5767_o[8];
  assign n6419_o = n5896_o[8];
  assign n6420_o = n5902_o[8];
  assign n6421_o = n5908_o[8];
  assign n6422_o = n6059_o[8];
  assign n6423_o = n6065_o[8];
  assign n6424_o = n6071_o[8];
  assign n6425_o = n6222_o[8];
  assign n6426_o = n6228_o[8];
  assign n6427_o = n6231_o[8];
  assign n6428_o = n6275_o[8];
  assign n6429_o = n5706_o[8];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = 1'b0;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6427_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6426_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6425_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6424_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6423_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6422_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6430_o = n6421_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6430_o = n6420_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6430_o = n6419_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6430_o = n6418_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6430_o = n6417_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6430_o = n6416_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6430_o = n6415_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6430_o = 1'b1;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6430_o = n6429_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6430_o = n6429_o;
      default: n6430_o = n6428_o;
    endcase
  assign n6431_o = n5750_o[9];
  assign n6432_o = n5755_o[9];
  assign n6433_o = n5760_o[9];
  assign n6434_o = n5767_o[9];
  assign n6435_o = n5896_o[9];
  assign n6436_o = n5902_o[9];
  assign n6437_o = n5908_o[9];
  assign n6438_o = n6059_o[9];
  assign n6439_o = n6065_o[9];
  assign n6440_o = n6071_o[9];
  assign n6441_o = n6222_o[9];
  assign n6442_o = n6228_o[9];
  assign n6443_o = n6231_o[9];
  assign n6444_o = n6275_o[9];
  assign n6445_o = n5706_o[9];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = 1'b0;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6443_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6442_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6441_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6440_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6439_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6438_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6446_o = n6437_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6446_o = n6436_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6446_o = n6435_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6446_o = n6434_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6446_o = n6433_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6446_o = n6432_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6446_o = n6431_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6446_o = n6445_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6446_o = n6445_o;
      default: n6446_o = n6444_o;
    endcase
  assign n6447_o = n5750_o[10];
  assign n6448_o = n5755_o[10];
  assign n6449_o = n5760_o[10];
  assign n6450_o = n5767_o[10];
  assign n6451_o = n5896_o[10];
  assign n6452_o = n5902_o[10];
  assign n6453_o = n5908_o[10];
  assign n6454_o = n6059_o[10];
  assign n6455_o = n6065_o[10];
  assign n6456_o = n6071_o[10];
  assign n6457_o = n6222_o[10];
  assign n6458_o = n6228_o[10];
  assign n6459_o = n6231_o[10];
  assign n6460_o = n6275_o[10];
  assign n6461_o = n5706_o[10];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = 1'b0;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6459_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6458_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6457_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6456_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6455_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6454_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6462_o = n6453_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6462_o = n6452_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6462_o = n6451_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6462_o = n6450_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6462_o = n6449_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6462_o = n6448_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6462_o = n6447_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6462_o = n6461_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6462_o = n6461_o;
      default: n6462_o = n6460_o;
    endcase
  assign n6463_o = n5717_o[0];
  assign n6464_o = n5750_o[11];
  assign n6465_o = n5755_o[11];
  assign n6466_o = n5760_o[11];
  assign n6467_o = n5767_o[11];
  assign n6468_o = n5896_o[11];
  assign n6469_o = n5902_o[11];
  assign n6470_o = n5908_o[11];
  assign n6471_o = n6059_o[11];
  assign n6472_o = n6065_o[11];
  assign n6473_o = n6071_o[11];
  assign n6474_o = n6222_o[11];
  assign n6475_o = n6228_o[11];
  assign n6476_o = n6231_o[11];
  assign n6477_o = n6275_o[11];
  assign n6478_o = n5706_o[11];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = 1'b0;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6476_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6475_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6474_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6473_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6472_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6471_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6479_o = n6470_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6479_o = n6469_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6479_o = n6468_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6479_o = n5772_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6479_o = n6467_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6479_o = n6466_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6479_o = n6465_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6479_o = n6464_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6479_o = n5744_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6479_o = n6463_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6479_o = n6478_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6479_o = n6478_o;
      default: n6479_o = n6477_o;
    endcase
  assign n6480_o = n5717_o[1];
  assign n6481_o = n5750_o[12];
  assign n6482_o = n5755_o[12];
  assign n6483_o = n5760_o[12];
  assign n6484_o = n5767_o[12];
  assign n6485_o = n5896_o[12];
  assign n6486_o = n5902_o[12];
  assign n6487_o = n5908_o[12];
  assign n6488_o = n6059_o[12];
  assign n6489_o = n6065_o[12];
  assign n6490_o = n6071_o[12];
  assign n6491_o = n6222_o[12];
  assign n6492_o = n6228_o[12];
  assign n6493_o = n6231_o[12];
  assign n6494_o = n6275_o[12];
  assign n6495_o = n5706_o[12];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6493_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6492_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6491_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6490_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6489_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6488_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6496_o = n6487_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6496_o = n6486_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6496_o = n6485_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6496_o = n6484_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6496_o = n6483_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6496_o = n6482_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6496_o = n6481_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6496_o = 1'b1;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6496_o = n6480_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6496_o = n6495_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6496_o = n6495_o;
      default: n6496_o = n6494_o;
    endcase
  assign n6497_o = n5750_o[15:13];
  assign n6498_o = n5755_o[15:13];
  assign n6499_o = n5760_o[15:13];
  assign n6500_o = n5767_o[15:13];
  assign n6501_o = n5896_o[15:13];
  assign n6502_o = n5902_o[15:13];
  assign n6503_o = n5908_o[15:13];
  assign n6504_o = n6059_o[15:13];
  assign n6505_o = n6065_o[15:13];
  assign n6506_o = n6071_o[15:13];
  assign n6507_o = n6222_o[15:13];
  assign n6508_o = n6228_o[15:13];
  assign n6509_o = n6231_o[15:13];
  assign n6510_o = n6275_o[15:13];
  assign n6511_o = n5706_o[15:13];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6509_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6508_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6507_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6506_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6505_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6504_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6512_o = n6503_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6512_o = n6502_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6512_o = n6501_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6512_o = n6500_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6512_o = n6499_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6512_o = n6498_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6512_o = n6497_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6512_o = n6511_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6512_o = n6511_o;
      default: n6512_o = n6510_o;
    endcase
  assign n6513_o = n5745_o[0];
  assign n6514_o = n5750_o[16];
  assign n6515_o = n5755_o[16];
  assign n6516_o = n5760_o[16];
  assign n6517_o = n5767_o[16];
  assign n6518_o = n5773_o[0];
  assign n6519_o = n5896_o[16];
  assign n6520_o = n5902_o[16];
  assign n6521_o = n5908_o[16];
  assign n6522_o = n6059_o[16];
  assign n6523_o = n6065_o[16];
  assign n6524_o = n6071_o[16];
  assign n6525_o = n6222_o[16];
  assign n6526_o = n6228_o[16];
  assign n6527_o = n6231_o[16];
  assign n6528_o = n6275_o[16];
  assign n6529_o = n5706_o[16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6527_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6526_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6525_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6524_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6523_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6522_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6530_o = n6521_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6530_o = n6520_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6530_o = n6519_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6530_o = n6518_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6530_o = n6517_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6530_o = n6516_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6530_o = n6515_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6530_o = n6514_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6530_o = n6513_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6530_o = n6529_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6530_o = n6529_o;
      default: n6530_o = n6528_o;
    endcase
  assign n6531_o = n5745_o[1];
  assign n6532_o = n5750_o[17];
  assign n6533_o = n5755_o[17];
  assign n6534_o = n5760_o[17];
  assign n6535_o = n5767_o[17];
  assign n6536_o = n5773_o[1];
  assign n6537_o = n5896_o[17];
  assign n6538_o = n5902_o[17];
  assign n6539_o = n5908_o[17];
  assign n6540_o = n6059_o[17];
  assign n6541_o = n6065_o[17];
  assign n6542_o = n6071_o[17];
  assign n6543_o = n6222_o[17];
  assign n6544_o = n6228_o[17];
  assign n6545_o = n6231_o[17];
  assign n6546_o = n6275_o[17];
  assign n6547_o = n5706_o[17];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6545_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6544_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6543_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6542_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6541_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6540_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6548_o = n6539_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6548_o = n6538_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6548_o = n6537_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6548_o = n6536_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6548_o = n6535_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6548_o = n6534_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6548_o = n6533_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6548_o = n6532_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6548_o = n6531_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6548_o = n5718_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6548_o = n6547_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6548_o = n6547_o;
      default: n6548_o = n6546_o;
    endcase
  assign n6549_o = n5745_o[3:2];
  assign n6550_o = n5750_o[19:18];
  assign n6551_o = n5755_o[19:18];
  assign n6552_o = n5760_o[19:18];
  assign n6553_o = n5767_o[19:18];
  assign n6554_o = n5773_o[3:2];
  assign n6555_o = n5896_o[19:18];
  assign n6556_o = n5902_o[19:18];
  assign n6557_o = n5908_o[19:18];
  assign n6558_o = n6059_o[19:18];
  assign n6559_o = n6065_o[19:18];
  assign n6560_o = n6071_o[19:18];
  assign n6561_o = n6222_o[19:18];
  assign n6562_o = n6228_o[19:18];
  assign n6563_o = n6231_o[19:18];
  assign n6564_o = n6275_o[19:18];
  assign n6565_o = n5706_o[19:18];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6563_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6562_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6561_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6560_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6559_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6558_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6566_o = n6557_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6566_o = n6556_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6566_o = n6555_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6566_o = n6554_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6566_o = n6553_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6566_o = n6552_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6566_o = n6551_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6566_o = n6550_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6566_o = n6549_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6566_o = n6565_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6566_o = n6565_o;
      default: n6566_o = n6564_o;
    endcase
  assign n6567_o = n5745_o[4];
  assign n6568_o = n5750_o[20];
  assign n6569_o = n5755_o[20];
  assign n6570_o = n5760_o[20];
  assign n6571_o = n5767_o[20];
  assign n6572_o = n5773_o[4];
  assign n6573_o = n5896_o[20];
  assign n6574_o = n5902_o[20];
  assign n6575_o = n5908_o[20];
  assign n6576_o = n6059_o[20];
  assign n6577_o = n6065_o[20];
  assign n6578_o = n6071_o[20];
  assign n6579_o = n6222_o[20];
  assign n6580_o = n6228_o[20];
  assign n6581_o = n6231_o[20];
  assign n6582_o = n6275_o[20];
  assign n6583_o = n5706_o[20];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = 1'b0;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6581_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6580_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6579_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6578_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6577_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6576_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6584_o = n6575_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6584_o = n6574_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6584_o = n6573_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6584_o = n6572_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6584_o = n6571_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6584_o = n6570_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6584_o = n6569_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6584_o = n6568_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6584_o = n6567_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6584_o = 1'b0;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6584_o = n6583_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6584_o = n6583_o;
      default: n6584_o = n6582_o;
    endcase
  assign n6585_o = n5745_o[5];
  assign n6586_o = n5750_o[21];
  assign n6587_o = n5755_o[21];
  assign n6588_o = n5760_o[21];
  assign n6589_o = n5767_o[21];
  assign n6590_o = n5773_o[5];
  assign n6591_o = n5896_o[21];
  assign n6592_o = n5902_o[21];
  assign n6593_o = n5908_o[21];
  assign n6594_o = n6059_o[21];
  assign n6595_o = n6065_o[21];
  assign n6596_o = n6071_o[21];
  assign n6597_o = n6222_o[21];
  assign n6598_o = n6228_o[21];
  assign n6599_o = n6231_o[21];
  assign n6600_o = n6275_o[21];
  assign n6601_o = n5706_o[21];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6599_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6598_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6597_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6596_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6595_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6594_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6602_o = n6593_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6602_o = n6592_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6602_o = n6591_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6602_o = n6590_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6602_o = n6589_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6602_o = n6588_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6602_o = n6587_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6602_o = n6586_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6602_o = n6585_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6602_o = n5722_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6602_o = n6601_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6602_o = n6601_o;
      default: n6602_o = n6600_o;
    endcase
  assign n6603_o = n5745_o[6];
  assign n6604_o = n5750_o[22];
  assign n6605_o = n5755_o[22];
  assign n6606_o = n5760_o[22];
  assign n6607_o = n5767_o[22];
  assign n6608_o = n5773_o[6];
  assign n6609_o = n5896_o[22];
  assign n6610_o = n5902_o[22];
  assign n6611_o = n5908_o[22];
  assign n6612_o = n6059_o[22];
  assign n6613_o = n6065_o[22];
  assign n6614_o = n6071_o[22];
  assign n6615_o = n6222_o[22];
  assign n6616_o = n6228_o[22];
  assign n6617_o = n6231_o[22];
  assign n6618_o = n6275_o[22];
  assign n6619_o = n5706_o[22];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6617_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6616_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6615_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6614_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6613_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6612_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6620_o = n6611_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6620_o = n6610_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6620_o = n6609_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6620_o = n6608_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6620_o = n6607_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6620_o = n6606_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6620_o = n6605_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6620_o = n6604_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6620_o = n6603_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6620_o = n6619_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6620_o = n6619_o;
      default: n6620_o = n6618_o;
    endcase
  assign n6621_o = n5745_o[7];
  assign n6622_o = n5750_o[23];
  assign n6623_o = n5755_o[23];
  assign n6624_o = n5760_o[23];
  assign n6625_o = n5767_o[23];
  assign n6626_o = n5773_o[7];
  assign n6627_o = n5896_o[23];
  assign n6628_o = n5902_o[23];
  assign n6629_o = n5908_o[23];
  assign n6630_o = n6059_o[23];
  assign n6631_o = n6065_o[23];
  assign n6632_o = n6071_o[23];
  assign n6633_o = n6222_o[23];
  assign n6634_o = n6228_o[23];
  assign n6635_o = n6231_o[23];
  assign n6636_o = n6275_o[23];
  assign n6637_o = n5706_o[23];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6635_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6634_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6633_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6632_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6631_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6630_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6638_o = n6629_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6638_o = n6628_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6638_o = n6627_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6638_o = n6626_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6638_o = n6625_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6638_o = n6624_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6638_o = n6623_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6638_o = n6622_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6638_o = n6621_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6638_o = 1'b1;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6638_o = n6637_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6638_o = n6637_o;
      default: n6638_o = n6636_o;
    endcase
  assign n6639_o = n5745_o[13:8];
  assign n6640_o = n5750_o[29:24];
  assign n6641_o = n5755_o[29:24];
  assign n6642_o = n5760_o[29:24];
  assign n6643_o = n5767_o[29:24];
  assign n6644_o = n5773_o[13:8];
  assign n6645_o = n5896_o[29:24];
  assign n6646_o = n5902_o[29:24];
  assign n6647_o = n5908_o[29:24];
  assign n6648_o = n6059_o[29:24];
  assign n6649_o = n6065_o[29:24];
  assign n6650_o = n6071_o[29:24];
  assign n6651_o = n6222_o[29:24];
  assign n6652_o = n6228_o[29:24];
  assign n6653_o = n6231_o[29:24];
  assign n6654_o = n6275_o[29:24];
  assign n6655_o = n5706_o[29:24];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6653_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6652_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6651_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6650_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6649_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6648_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6656_o = n6647_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6656_o = n6646_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6656_o = n6645_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6656_o = n6644_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6656_o = n6643_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6656_o = n6642_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6656_o = n6641_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6656_o = n6640_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6656_o = n6639_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6656_o = n6655_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6656_o = n6655_o;
      default: n6656_o = n6654_o;
    endcase
  assign n6657_o = n5745_o[14];
  assign n6658_o = n5750_o[30];
  assign n6659_o = n5755_o[30];
  assign n6660_o = n5760_o[30];
  assign n6661_o = n5767_o[30];
  assign n6662_o = n5773_o[14];
  assign n6663_o = n5896_o[30];
  assign n6664_o = n5902_o[30];
  assign n6665_o = n5908_o[30];
  assign n6666_o = n6059_o[30];
  assign n6667_o = n6065_o[30];
  assign n6668_o = n6071_o[30];
  assign n6669_o = n6222_o[30];
  assign n6670_o = n6228_o[30];
  assign n6671_o = n6231_o[30];
  assign n6672_o = n6275_o[30];
  assign n6673_o = n5706_o[30];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = 1'b0;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6671_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6670_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6669_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6668_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6667_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6666_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6674_o = n6665_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6674_o = n6664_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6674_o = n6663_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6674_o = n6662_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6674_o = n6661_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6674_o = n6660_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6674_o = n6659_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6674_o = n6658_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6674_o = n6657_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6674_o = 1'b1;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6674_o = n6673_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6674_o = n6673_o;
      default: n6674_o = n6672_o;
    endcase
  assign n6675_o = n5745_o[15];
  assign n6676_o = n5750_o[31];
  assign n6677_o = n5755_o[31];
  assign n6678_o = n5760_o[31];
  assign n6679_o = n5767_o[31];
  assign n6680_o = n5773_o[15];
  assign n6681_o = n5896_o[31];
  assign n6682_o = n5902_o[31];
  assign n6683_o = n5908_o[31];
  assign n6684_o = n6059_o[31];
  assign n6685_o = n6065_o[31];
  assign n6686_o = n6071_o[31];
  assign n6687_o = n6222_o[31];
  assign n6688_o = n6228_o[31];
  assign n6689_o = n6231_o[31];
  assign n6690_o = n6275_o[31];
  assign n6691_o = n5706_o[31];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2126:7  */
  always @*
    case (n6276_o)
      120'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = 1'b0;
      120'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6689_o;
      120'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6688_o;
      120'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6687_o;
      120'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6686_o;
      120'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6685_o;
      120'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6684_o;
      120'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6692_o = n6683_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6692_o = n6682_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6692_o = n6681_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6692_o = n6680_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6692_o = n6679_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6692_o = n5763_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6692_o = n6678_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6692_o = n6677_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6692_o = n6676_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6692_o = n6675_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6692_o = 1'b0;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6692_o = n6691_o;
      120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6692_o = n6691_o;
      default: n6692_o = n6690_o;
    endcase
  assign n6716_o = {n6692_o, n6674_o, n6656_o, n6638_o, n6620_o, n6602_o, n6584_o, n6566_o, n6548_o, n6530_o, n6512_o, n6496_o, n6479_o, n6462_o, n6446_o, n6430_o, n6414_o, n6398_o, n6382_o, n6366_o, n6348_o, n6330_o, n6312_o, n6294_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2396:25  */
  assign n6722_o = csr[11:10];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2396:50  */
  assign n6723_o = csr[8];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2396:40  */
  assign n6724_o = {n6722_o, n6723_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2396:64  */
  assign n6725_o = csr[8];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2396:54  */
  assign n6726_o = {n6724_o, n6725_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2396:78  */
  assign n6727_o = csr[7:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2396:68  */
  assign n6728_o = {n6726_o, n6727_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2396:102  */
  assign n6729_o = csr[14];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2396:92  */
  assign n6730_o = n6729_o ? n6728_o : 12'b000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2399:22  */
  assign n6732_o = csr[79:48];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2414:13  */
  assign n6736_o = csr[12];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2414:36  */
  assign n6737_o = csr[11:8];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2414:50  */
  assign n6739_o = n6737_o == 4'b1011;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2414:23  */
  assign n6740_o = n6736_o & n6739_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2415:19  */
  assign n6741_o = csr[7];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2415:23  */
  assign n6742_o = ~n6741_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:47  */
  assign n6743_o = csr[4:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:47  */
  assign n6748_o = csr[4:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2415:7  */
  assign n6753_o = n6742_o ? n8562_o : 32'b00000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2415:7  */
  assign n6754_o = n6742_o ? 32'b00000000000000000000000000000000 : n8697_o;
  assign n6755_o = {n6754_o, n6753_o};
  assign n6756_o = {32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2414:5  */
  assign n6757_o = n6740_o ? n6755_o : n6756_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n6760_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n6765_o = cnt[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n6766_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n6767_o = cnt[3198:3167];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n6768_o = n6765_o ? n6766_o : n6767_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n6769_o = cnt[3199];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n6770_o = cnt[32];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n6771_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n6772_o = cnt[2143:2112];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n6773_o = cnt[3231];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n6774_o = {31'b0, n6773_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n6775_o = n6772_o + n6774_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n6776_o = n6770_o ? n6771_o : n6775_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n6787_o = cnt[1119:1088];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n6789_o = {1'b0, n6787_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n6791_o = n6789_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n6792_o = cnt[64];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n6793_o = n6792_o ? n6791_o : n6798_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n6794_o = cnt[1119:1088];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n6796_o = {1'b0, n6794_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n6798_o = n6796_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n6800_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n6805_o = cnt[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n6806_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n6807_o = cnt[3165:3134];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n6808_o = n6805_o ? n6806_o : n6807_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n6809_o = cnt[3166];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n6810_o = cnt[33];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n6811_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n6812_o = cnt[2111:2080];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n6813_o = cnt[3230];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n6814_o = {31'b0, n6813_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n6815_o = n6812_o + n6814_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n6816_o = n6810_o ? n6811_o : n6815_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n6827_o = cnt[1087:1056];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n6829_o = {1'b0, n6827_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n6831_o = n6829_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n6832_o = cnt[65];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n6833_o = n6832_o ? n6831_o : n6838_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n6834_o = cnt[1087:1056];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n6836_o = {1'b0, n6834_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n6838_o = n6836_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n6840_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n6845_o = cnt[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n6846_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n6847_o = cnt[3132:3101];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n6848_o = n6845_o ? n6846_o : n6847_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n6849_o = cnt[3133];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n6850_o = cnt[34];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n6851_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n6852_o = cnt[2079:2048];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n6853_o = cnt[3229];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n6854_o = {31'b0, n6853_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n6855_o = n6852_o + n6854_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n6856_o = n6850_o ? n6851_o : n6855_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n6867_o = cnt[1055:1024];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n6869_o = {1'b0, n6867_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n6871_o = n6869_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n6872_o = cnt[66];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n6873_o = n6872_o ? n6871_o : n6878_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n6874_o = cnt[1055:1024];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n6876_o = {1'b0, n6874_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n6878_o = n6876_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n6880_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n6885_o = cnt[3];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n6886_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n6887_o = cnt[3099:3068];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n6888_o = n6885_o ? n6886_o : n6887_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n6889_o = cnt[3100];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n6890_o = cnt[35];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n6891_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n6892_o = cnt[2047:2016];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n6893_o = cnt[3228];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n6894_o = {31'b0, n6893_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n6895_o = n6892_o + n6894_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n6896_o = n6890_o ? n6891_o : n6895_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n6907_o = cnt[1023:992];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n6909_o = {1'b0, n6907_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n6911_o = n6909_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n6912_o = cnt[67];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n6913_o = n6912_o ? n6911_o : n6918_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n6914_o = cnt[1023:992];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n6916_o = {1'b0, n6914_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n6918_o = n6916_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n6920_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n6925_o = cnt[4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n6926_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n6927_o = cnt[3066:3035];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n6928_o = n6925_o ? n6926_o : n6927_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n6929_o = cnt[3067];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n6930_o = cnt[36];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n6931_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n6932_o = cnt[2015:1984];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n6933_o = cnt[3227];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n6934_o = {31'b0, n6933_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n6935_o = n6932_o + n6934_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n6936_o = n6930_o ? n6931_o : n6935_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n6947_o = cnt[991:960];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n6949_o = {1'b0, n6947_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n6951_o = n6949_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n6952_o = cnt[68];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n6953_o = n6952_o ? n6951_o : n6958_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n6954_o = cnt[991:960];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n6956_o = {1'b0, n6954_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n6958_o = n6956_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n6960_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n6965_o = cnt[5];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n6966_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n6967_o = cnt[3033:3002];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n6968_o = n6965_o ? n6966_o : n6967_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n6969_o = cnt[3034];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n6970_o = cnt[37];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n6971_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n6972_o = cnt[1983:1952];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n6973_o = cnt[3226];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n6974_o = {31'b0, n6973_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n6975_o = n6972_o + n6974_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n6976_o = n6970_o ? n6971_o : n6975_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n6987_o = cnt[959:928];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n6989_o = {1'b0, n6987_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n6991_o = n6989_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n6992_o = cnt[69];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n6993_o = n6992_o ? n6991_o : n6998_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n6994_o = cnt[959:928];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n6996_o = {1'b0, n6994_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n6998_o = n6996_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7000_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7005_o = cnt[6];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7006_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7007_o = cnt[3000:2969];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7008_o = n7005_o ? n7006_o : n7007_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7009_o = cnt[3001];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7010_o = cnt[38];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7011_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7012_o = cnt[1951:1920];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7013_o = cnt[3225];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7014_o = {31'b0, n7013_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7015_o = n7012_o + n7014_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7016_o = n7010_o ? n7011_o : n7015_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7027_o = cnt[927:896];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7029_o = {1'b0, n7027_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7031_o = n7029_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7032_o = cnt[70];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7033_o = n7032_o ? n7031_o : n7038_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7034_o = cnt[927:896];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7036_o = {1'b0, n7034_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7038_o = n7036_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7040_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7045_o = cnt[7];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7046_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7047_o = cnt[2967:2936];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7048_o = n7045_o ? n7046_o : n7047_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7049_o = cnt[2968];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7050_o = cnt[39];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7051_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7052_o = cnt[1919:1888];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7053_o = cnt[3224];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7054_o = {31'b0, n7053_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7055_o = n7052_o + n7054_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7056_o = n7050_o ? n7051_o : n7055_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7067_o = cnt[895:864];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7069_o = {1'b0, n7067_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7071_o = n7069_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7072_o = cnt[71];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7073_o = n7072_o ? n7071_o : n7078_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7074_o = cnt[895:864];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7076_o = {1'b0, n7074_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7078_o = n7076_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7080_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7085_o = cnt[8];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7086_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7087_o = cnt[2934:2903];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7088_o = n7085_o ? n7086_o : n7087_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7089_o = cnt[2935];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7090_o = cnt[40];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7091_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7092_o = cnt[1887:1856];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7093_o = cnt[3223];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7094_o = {31'b0, n7093_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7095_o = n7092_o + n7094_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7096_o = n7090_o ? n7091_o : n7095_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7107_o = cnt[863:832];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7109_o = {1'b0, n7107_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7111_o = n7109_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7112_o = cnt[72];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7113_o = n7112_o ? n7111_o : n7118_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7114_o = cnt[863:832];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7116_o = {1'b0, n7114_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7118_o = n7116_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7120_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7125_o = cnt[9];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7126_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7127_o = cnt[2901:2870];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7128_o = n7125_o ? n7126_o : n7127_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7129_o = cnt[2902];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7130_o = cnt[41];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7131_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7132_o = cnt[1855:1824];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7133_o = cnt[3222];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7134_o = {31'b0, n7133_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7135_o = n7132_o + n7134_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7136_o = n7130_o ? n7131_o : n7135_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7147_o = cnt[831:800];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7149_o = {1'b0, n7147_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7151_o = n7149_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7152_o = cnt[73];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7153_o = n7152_o ? n7151_o : n7158_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7154_o = cnt[831:800];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7156_o = {1'b0, n7154_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7158_o = n7156_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7160_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7165_o = cnt[10];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7166_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7167_o = cnt[2868:2837];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7168_o = n7165_o ? n7166_o : n7167_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7169_o = cnt[2869];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7170_o = cnt[42];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7171_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7172_o = cnt[1823:1792];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7173_o = cnt[3221];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7174_o = {31'b0, n7173_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7175_o = n7172_o + n7174_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7176_o = n7170_o ? n7171_o : n7175_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7187_o = cnt[799:768];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7189_o = {1'b0, n7187_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7191_o = n7189_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7192_o = cnt[74];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7193_o = n7192_o ? n7191_o : n7198_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7194_o = cnt[799:768];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7196_o = {1'b0, n7194_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7198_o = n7196_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7200_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7205_o = cnt[11];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7206_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7207_o = cnt[2835:2804];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7208_o = n7205_o ? n7206_o : n7207_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7209_o = cnt[2836];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7210_o = cnt[43];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7211_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7212_o = cnt[1791:1760];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7213_o = cnt[3220];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7214_o = {31'b0, n7213_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7215_o = n7212_o + n7214_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7216_o = n7210_o ? n7211_o : n7215_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7227_o = cnt[767:736];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7229_o = {1'b0, n7227_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7231_o = n7229_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7232_o = cnt[75];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7233_o = n7232_o ? n7231_o : n7238_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7234_o = cnt[767:736];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7236_o = {1'b0, n7234_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7238_o = n7236_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7240_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7245_o = cnt[12];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7246_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7247_o = cnt[2802:2771];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7248_o = n7245_o ? n7246_o : n7247_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7249_o = cnt[2803];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7250_o = cnt[44];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7251_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7252_o = cnt[1759:1728];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7253_o = cnt[3219];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7254_o = {31'b0, n7253_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7255_o = n7252_o + n7254_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7256_o = n7250_o ? n7251_o : n7255_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7267_o = cnt[735:704];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7269_o = {1'b0, n7267_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7271_o = n7269_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7272_o = cnt[76];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7273_o = n7272_o ? n7271_o : n7278_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7274_o = cnt[735:704];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7276_o = {1'b0, n7274_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7278_o = n7276_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7280_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7285_o = cnt[13];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7286_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7287_o = cnt[2769:2738];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7288_o = n7285_o ? n7286_o : n7287_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7289_o = cnt[2770];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7290_o = cnt[45];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7291_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7292_o = cnt[1727:1696];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7293_o = cnt[3218];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7294_o = {31'b0, n7293_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7295_o = n7292_o + n7294_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7296_o = n7290_o ? n7291_o : n7295_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7307_o = cnt[703:672];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7309_o = {1'b0, n7307_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7311_o = n7309_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7312_o = cnt[77];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7313_o = n7312_o ? n7311_o : n7318_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7314_o = cnt[703:672];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7316_o = {1'b0, n7314_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7318_o = n7316_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7320_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7325_o = cnt[14];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7326_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7327_o = cnt[2736:2705];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7328_o = n7325_o ? n7326_o : n7327_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7329_o = cnt[2737];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7330_o = cnt[46];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7331_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7332_o = cnt[1695:1664];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7333_o = cnt[3217];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7334_o = {31'b0, n7333_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7335_o = n7332_o + n7334_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7336_o = n7330_o ? n7331_o : n7335_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7347_o = cnt[671:640];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7349_o = {1'b0, n7347_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7351_o = n7349_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7352_o = cnt[78];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7353_o = n7352_o ? n7351_o : n7358_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7354_o = cnt[671:640];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7356_o = {1'b0, n7354_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7358_o = n7356_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7360_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7365_o = cnt[15];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7366_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7367_o = cnt[2703:2672];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7368_o = n7365_o ? n7366_o : n7367_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7369_o = cnt[2704];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7370_o = cnt[47];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7371_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7372_o = cnt[1663:1632];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7373_o = cnt[3216];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7374_o = {31'b0, n7373_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7375_o = n7372_o + n7374_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7376_o = n7370_o ? n7371_o : n7375_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7387_o = cnt[639:608];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7389_o = {1'b0, n7387_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7391_o = n7389_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7392_o = cnt[79];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7393_o = n7392_o ? n7391_o : n7398_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7394_o = cnt[639:608];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7396_o = {1'b0, n7394_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7398_o = n7396_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7400_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7405_o = cnt[16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7406_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7407_o = cnt[2670:2639];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7408_o = n7405_o ? n7406_o : n7407_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7409_o = cnt[2671];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7410_o = cnt[48];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7411_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7412_o = cnt[1631:1600];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7413_o = cnt[3215];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7414_o = {31'b0, n7413_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7415_o = n7412_o + n7414_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7416_o = n7410_o ? n7411_o : n7415_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7427_o = cnt[607:576];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7429_o = {1'b0, n7427_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7431_o = n7429_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7432_o = cnt[80];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7433_o = n7432_o ? n7431_o : n7438_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7434_o = cnt[607:576];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7436_o = {1'b0, n7434_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7438_o = n7436_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7440_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7445_o = cnt[17];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7446_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7447_o = cnt[2637:2606];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7448_o = n7445_o ? n7446_o : n7447_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7449_o = cnt[2638];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7450_o = cnt[49];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7451_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7452_o = cnt[1599:1568];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7453_o = cnt[3214];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7454_o = {31'b0, n7453_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7455_o = n7452_o + n7454_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7456_o = n7450_o ? n7451_o : n7455_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7467_o = cnt[575:544];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7469_o = {1'b0, n7467_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7471_o = n7469_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7472_o = cnt[81];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7473_o = n7472_o ? n7471_o : n7478_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7474_o = cnt[575:544];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7476_o = {1'b0, n7474_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7478_o = n7476_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7480_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7485_o = cnt[18];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7486_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7487_o = cnt[2604:2573];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7488_o = n7485_o ? n7486_o : n7487_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7489_o = cnt[2605];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7490_o = cnt[50];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7491_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7492_o = cnt[1567:1536];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7493_o = cnt[3213];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7494_o = {31'b0, n7493_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7495_o = n7492_o + n7494_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7496_o = n7490_o ? n7491_o : n7495_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7507_o = cnt[543:512];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7509_o = {1'b0, n7507_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7511_o = n7509_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7512_o = cnt[82];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7513_o = n7512_o ? n7511_o : n7518_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7514_o = cnt[543:512];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7516_o = {1'b0, n7514_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7518_o = n7516_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7520_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7525_o = cnt[19];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7526_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7527_o = cnt[2571:2540];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7528_o = n7525_o ? n7526_o : n7527_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7529_o = cnt[2572];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7530_o = cnt[51];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7531_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7532_o = cnt[1535:1504];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7533_o = cnt[3212];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7534_o = {31'b0, n7533_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7535_o = n7532_o + n7534_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7536_o = n7530_o ? n7531_o : n7535_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7547_o = cnt[511:480];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7549_o = {1'b0, n7547_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7551_o = n7549_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7552_o = cnt[83];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7553_o = n7552_o ? n7551_o : n7558_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7554_o = cnt[511:480];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7556_o = {1'b0, n7554_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7558_o = n7556_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7560_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7565_o = cnt[20];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7566_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7567_o = cnt[2538:2507];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7568_o = n7565_o ? n7566_o : n7567_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7569_o = cnt[2539];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7570_o = cnt[52];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7571_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7572_o = cnt[1503:1472];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7573_o = cnt[3211];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7574_o = {31'b0, n7573_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7575_o = n7572_o + n7574_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7576_o = n7570_o ? n7571_o : n7575_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7587_o = cnt[479:448];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7589_o = {1'b0, n7587_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7591_o = n7589_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7592_o = cnt[84];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7593_o = n7592_o ? n7591_o : n7598_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7594_o = cnt[479:448];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7596_o = {1'b0, n7594_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7598_o = n7596_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7600_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7605_o = cnt[21];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7606_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7607_o = cnt[2505:2474];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7608_o = n7605_o ? n7606_o : n7607_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7609_o = cnt[2506];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7610_o = cnt[53];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7611_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7612_o = cnt[1471:1440];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7613_o = cnt[3210];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7614_o = {31'b0, n7613_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7615_o = n7612_o + n7614_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7616_o = n7610_o ? n7611_o : n7615_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7627_o = cnt[447:416];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7629_o = {1'b0, n7627_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7631_o = n7629_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7632_o = cnt[85];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7633_o = n7632_o ? n7631_o : n7638_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7634_o = cnt[447:416];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7636_o = {1'b0, n7634_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7638_o = n7636_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7640_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7645_o = cnt[22];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7646_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7647_o = cnt[2472:2441];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7648_o = n7645_o ? n7646_o : n7647_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7649_o = cnt[2473];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7650_o = cnt[54];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7651_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7652_o = cnt[1439:1408];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7653_o = cnt[3209];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7654_o = {31'b0, n7653_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7655_o = n7652_o + n7654_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7656_o = n7650_o ? n7651_o : n7655_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7667_o = cnt[415:384];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7669_o = {1'b0, n7667_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7671_o = n7669_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7672_o = cnt[86];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7673_o = n7672_o ? n7671_o : n7678_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7674_o = cnt[415:384];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7676_o = {1'b0, n7674_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7678_o = n7676_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7680_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7685_o = cnt[23];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7686_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7687_o = cnt[2439:2408];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7688_o = n7685_o ? n7686_o : n7687_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7689_o = cnt[2440];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7690_o = cnt[55];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7691_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7692_o = cnt[1407:1376];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7693_o = cnt[3208];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7694_o = {31'b0, n7693_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7695_o = n7692_o + n7694_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7696_o = n7690_o ? n7691_o : n7695_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7707_o = cnt[383:352];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7709_o = {1'b0, n7707_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7711_o = n7709_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7712_o = cnt[87];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7713_o = n7712_o ? n7711_o : n7718_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7714_o = cnt[383:352];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7716_o = {1'b0, n7714_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7718_o = n7716_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7720_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7725_o = cnt[24];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7726_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7727_o = cnt[2406:2375];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7728_o = n7725_o ? n7726_o : n7727_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7729_o = cnt[2407];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7730_o = cnt[56];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7731_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7732_o = cnt[1375:1344];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7733_o = cnt[3207];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7734_o = {31'b0, n7733_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7735_o = n7732_o + n7734_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7736_o = n7730_o ? n7731_o : n7735_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7747_o = cnt[351:320];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7749_o = {1'b0, n7747_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7751_o = n7749_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7752_o = cnt[88];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7753_o = n7752_o ? n7751_o : n7758_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7754_o = cnt[351:320];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7756_o = {1'b0, n7754_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7758_o = n7756_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7760_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7765_o = cnt[25];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7766_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7767_o = cnt[2373:2342];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7768_o = n7765_o ? n7766_o : n7767_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7769_o = cnt[2374];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7770_o = cnt[57];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7771_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7772_o = cnt[1343:1312];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7773_o = cnt[3206];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7774_o = {31'b0, n7773_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7775_o = n7772_o + n7774_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7776_o = n7770_o ? n7771_o : n7775_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7787_o = cnt[319:288];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7789_o = {1'b0, n7787_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7791_o = n7789_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7792_o = cnt[89];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7793_o = n7792_o ? n7791_o : n7798_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7794_o = cnt[319:288];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7796_o = {1'b0, n7794_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7798_o = n7796_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7800_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7805_o = cnt[26];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7806_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7807_o = cnt[2340:2309];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7808_o = n7805_o ? n7806_o : n7807_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7809_o = cnt[2341];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7810_o = cnt[58];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7811_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7812_o = cnt[1311:1280];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7813_o = cnt[3205];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7814_o = {31'b0, n7813_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7815_o = n7812_o + n7814_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7816_o = n7810_o ? n7811_o : n7815_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7827_o = cnt[287:256];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7829_o = {1'b0, n7827_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7831_o = n7829_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7832_o = cnt[90];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7833_o = n7832_o ? n7831_o : n7838_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7834_o = cnt[287:256];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7836_o = {1'b0, n7834_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7838_o = n7836_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7840_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7845_o = cnt[27];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7846_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7847_o = cnt[2307:2276];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7848_o = n7845_o ? n7846_o : n7847_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7849_o = cnt[2308];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7850_o = cnt[59];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7851_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7852_o = cnt[1279:1248];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7853_o = cnt[3204];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7854_o = {31'b0, n7853_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7855_o = n7852_o + n7854_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7856_o = n7850_o ? n7851_o : n7855_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7867_o = cnt[255:224];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7869_o = {1'b0, n7867_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7871_o = n7869_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7872_o = cnt[91];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7873_o = n7872_o ? n7871_o : n7878_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7874_o = cnt[255:224];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7876_o = {1'b0, n7874_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7878_o = n7876_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7880_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7885_o = cnt[28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7886_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7887_o = cnt[2274:2243];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7888_o = n7885_o ? n7886_o : n7887_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7889_o = cnt[2275];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7890_o = cnt[60];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7891_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7892_o = cnt[1247:1216];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7893_o = cnt[3203];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7894_o = {31'b0, n7893_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7895_o = n7892_o + n7894_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7896_o = n7890_o ? n7891_o : n7895_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7907_o = cnt[223:192];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7909_o = {1'b0, n7907_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7911_o = n7909_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7912_o = cnt[92];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7913_o = n7912_o ? n7911_o : n7918_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7914_o = cnt[223:192];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7916_o = {1'b0, n7914_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7918_o = n7916_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7920_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7925_o = cnt[29];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7926_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7927_o = cnt[2241:2210];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7928_o = n7925_o ? n7926_o : n7927_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7929_o = cnt[2242];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7930_o = cnt[61];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7931_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7932_o = cnt[1215:1184];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7933_o = cnt[3202];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7934_o = {31'b0, n7933_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7935_o = n7932_o + n7934_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7936_o = n7930_o ? n7931_o : n7935_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7947_o = cnt[191:160];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7949_o = {1'b0, n7947_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7951_o = n7949_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7952_o = cnt[93];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7953_o = n7952_o ? n7951_o : n7958_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7954_o = cnt[191:160];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7956_o = {1'b0, n7954_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7958_o = n7956_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n7960_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n7965_o = cnt[30];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n7966_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n7967_o = cnt[2208:2177];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n7968_o = n7965_o ? n7966_o : n7967_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n7969_o = cnt[2209];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n7970_o = cnt[62];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n7971_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n7972_o = cnt[1183:1152];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n7973_o = cnt[3201];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7974_o = {31'b0, n7973_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n7975_o = n7972_o + n7974_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n7976_o = n7970_o ? n7971_o : n7975_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n7987_o = cnt[159:128];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n7989_o = {1'b0, n7987_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n7991_o = n7989_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n7992_o = cnt[94];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n7993_o = n7992_o ? n7991_o : n7998_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n7994_o = cnt[159:128];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n7996_o = {1'b0, n7994_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n7998_o = n7996_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:18  */
  assign n8000_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:22  */
  assign n8005_o = cnt[31];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2436:28  */
  assign n8006_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2438:34  */
  assign n8007_o = cnt[2175:2144];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2435:9  */
  assign n8008_o = n8005_o ? n8006_o : n8007_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2440:36  */
  assign n8009_o = cnt[2176];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:22  */
  assign n8010_o = cnt[63];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2443:28  */
  assign n8011_o = csr[47:16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:57  */
  assign n8012_o = cnt[1151:1120];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:80  */
  assign n8013_o = cnt[3200];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n8014_o = {31'b0, n8013_o};  //  uext
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2445:62  */
  assign n8015_o = n8012_o + n8014_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2442:9  */
  assign n8016_o = n8010_o ? n8011_o : n8015_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:58  */
  assign n8027_o = cnt[127:96];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:50  */
  assign n8029_o = {1'b0, n8027_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:63  */
  assign n8031_o = n8029_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:81  */
  assign n8032_o = cnt[95];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2451:68  */
  assign n8033_o = n8032_o ? n8031_o : n8038_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:58  */
  assign n8034_o = cnt[127:96];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:50  */
  assign n8036_o = {1'b0, n8034_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2452:63  */
  assign n8038_o = n8036_o + 33'b000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2462:29  */
  assign n8040_o = cnt[1119:1088];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2463:29  */
  assign n8043_o = cnt[2143:2112];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2464:29  */
  assign n8046_o = cnt[1119:1088];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2465:29  */
  assign n8048_o = cnt[2143:2112];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2466:29  */
  assign n8050_o = cnt[1055:1024];
  assign n8051_o = n8041_o[927:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2467:29  */
  assign n8052_o = cnt[2079:2048];
  assign n8053_o = n8044_o[927:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2491:30  */
  assign n8058_o = cnt_event[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2491:76  */
  assign n8059_o = csr[288];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2491:55  */
  assign n8060_o = ~n8059_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2491:50  */
  assign n8061_o = n8058_o & n8060_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2491:101  */
  assign n8062_o = debug_ctrl[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2491:86  */
  assign n8063_o = ~n8062_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2491:81  */
  assign n8064_o = n8061_o & n8063_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2492:30  */
  assign n8066_o = cnt_event[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2492:76  */
  assign n8067_o = csr[289];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2492:55  */
  assign n8068_o = ~n8067_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2492:50  */
  assign n8069_o = n8066_o & n8068_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2492:101  */
  assign n8070_o = debug_ctrl[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2492:86  */
  assign n8071_o = ~n8070_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2492:81  */
  assign n8072_o = n8069_o & n8071_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2493:30  */
  assign n8074_o = cnt_event[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2493:76  */
  assign n8075_o = csr[290];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2493:55  */
  assign n8076_o = ~n8075_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2493:50  */
  assign n8077_o = n8074_o & n8076_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2493:101  */
  assign n8078_o = debug_ctrl[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2493:86  */
  assign n8079_o = ~n8078_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2493:81  */
  assign n8080_o = n8077_o & n8079_o;
  assign n8081_o = n8057_o[31:3];
  assign n8082_o = {n8081_o, n8080_o, n8072_o, n8064_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2502:65  */
  assign n8087_o = execute_engine[215];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2502:71  */
  assign n8088_o = ~n8087_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2502:44  */
  assign n8089_o = n8088_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2504:65  */
  assign n8093_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2504:71  */
  assign n8095_o = n8093_o == 4'b0101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2504:44  */
  assign n8096_o = n8095_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2507:65  */
  assign n8099_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2507:71  */
  assign n8101_o = n8099_o == 4'b0101;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2507:105  */
  assign n8102_o = execute_engine[80];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2507:85  */
  assign n8103_o = n8101_o & n8102_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2507:44  */
  assign n8104_o = n8103_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2508:63  */
  assign n8107_o = fetch_engine[1:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2508:71  */
  assign n8109_o = n8107_o == 2'b10;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2508:103  */
  assign n8110_o = fetch_engine[3:2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2508:116  */
  assign n8112_o = n8110_o == 2'b10;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2508:85  */
  assign n8113_o = n8109_o & n8112_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2508:44  */
  assign n8114_o = n8113_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2509:65  */
  assign n8117_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2509:71  */
  assign n8119_o = n8117_o == 4'b0001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2509:105  */
  assign n8120_o = execute_engine[11:8];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2509:116  */
  assign n8122_o = n8120_o == 4'b0001;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2509:85  */
  assign n8123_o = n8119_o & n8122_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2509:44  */
  assign n8124_o = n8123_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2510:65  */
  assign n8127_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2510:71  */
  assign n8129_o = n8127_o == 4'b0110;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2510:44  */
  assign n8130_o = n8129_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2512:55  */
  assign n8133_o = ctrl[39];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2512:108  */
  assign n8134_o = execute_engine[21];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2512:131  */
  assign n8135_o = ~n8134_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2512:83  */
  assign n8136_o = n8133_o & n8135_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2512:44  */
  assign n8137_o = n8136_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2513:55  */
  assign n8140_o = ctrl[39];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2513:108  */
  assign n8141_o = execute_engine[21];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2513:83  */
  assign n8142_o = n8140_o & n8141_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2513:44  */
  assign n8143_o = n8142_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2514:65  */
  assign n8146_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2514:71  */
  assign n8148_o = n8146_o == 4'b1010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2514:103  */
  assign n8149_o = execute_engine[15:12];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2514:115  */
  assign n8151_o = n8149_o == 4'b1010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2514:83  */
  assign n8152_o = n8148_o & n8151_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2514:44  */
  assign n8153_o = n8152_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2516:65  */
  assign n8156_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2516:71  */
  assign n8158_o = n8156_o == 4'b0111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2516:108  */
  assign n8159_o = execute_engine[18];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2516:83  */
  assign n8160_o = n8158_o & n8159_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2516:44  */
  assign n8161_o = n8160_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2517:65  */
  assign n8164_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2517:71  */
  assign n8166_o = n8164_o == 4'b0111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2517:108  */
  assign n8167_o = execute_engine[18];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2517:131  */
  assign n8168_o = ~n8167_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2517:83  */
  assign n8169_o = n8166_o & n8168_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2517:44  */
  assign n8170_o = n8169_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2518:65  */
  assign n8173_o = execute_engine[3:0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2518:71  */
  assign n8175_o = n8173_o == 4'b0000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2518:103  */
  assign n8176_o = execute_engine[11:8];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2518:114  */
  assign n8178_o = n8176_o == 4'b0111;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2518:83  */
  assign n8179_o = n8175_o & n8178_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2519:108  */
  assign n8180_o = execute_engine[18];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2519:131  */
  assign n8181_o = ~n8180_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2518:124  */
  assign n8182_o = n8179_o & n8181_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2518:44  */
  assign n8183_o = n8182_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2521:60  */
  assign n8186_o = trap_ctrl[95];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2521:44  */
  assign n8187_o = n8186_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2522:60  */
  assign n8190_o = trap_ctrl[95];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2522:96  */
  assign n8191_o = trap_ctrl[61:55];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2522:102  */
  assign n8193_o = n8191_o == 7'b0000010;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2522:81  */
  assign n8194_o = n8190_o & n8193_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2522:44  */
  assign n8195_o = n8194_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2533:16  */
  assign n8198_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2568:29  */
  assign n8213_o = 1'b1 ? 1'b0 : 1'b1;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2571:64  */
  assign n8215_o = debug_ctrl[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2571:49  */
  assign n8216_o = ~n8215_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2571:44  */
  assign n8217_o = hw_trigger_fire & n8216_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2571:81  */
  assign n8218_o = csr[432];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2571:73  */
  assign n8219_o = n8217_o & n8218_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2571:103  */
  assign n8220_o = csr[433];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2571:95  */
  assign n8221_o = n8219_o & n8220_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2572:38  */
  assign n8222_o = trap_ctrl[101];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2572:66  */
  assign n8223_o = debug_ctrl[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2573:38  */
  assign n8224_o = csr[120];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2573:57  */
  assign n8225_o = csr[328];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2573:49  */
  assign n8226_o = n8224_o & n8225_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2572:74  */
  assign n8227_o = n8223_o | n8226_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2574:38  */
  assign n8228_o = csr[120];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2574:30  */
  assign n8229_o = ~n8228_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2574:57  */
  assign n8230_o = csr[329];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2574:49  */
  assign n8231_o = n8229_o & n8230_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2573:71  */
  assign n8232_o = n8227_o | n8231_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2572:50  */
  assign n8233_o = n8222_o & n8232_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2575:39  */
  assign n8234_o = debug_ctrl[8];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2575:72  */
  assign n8235_o = debug_ctrl[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2575:57  */
  assign n8236_o = ~n8235_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2575:52  */
  assign n8237_o = n8234_o & n8236_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2576:32  */
  assign n8238_o = csr[330];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2576:62  */
  assign n8239_o = debug_ctrl[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2576:47  */
  assign n8240_o = ~n8239_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2576:42  */
  assign n8241_o = n8238_o & n8240_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2583:36  */
  assign n8244_o = csr[328];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2586:36  */
  assign n8247_o = csr[329];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2586:49  */
  assign n8249_o = 1'b0 ? n8247_o : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2590:36  */
  assign n8254_o = csr[334:332];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2594:36  */
  assign n8258_o = csr[330];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2595:47  */
  assign n8259_o = csr[331];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2595:47  */
  assign n8260_o = csr[331];
  assign n8261_o = {n8259_o, n8260_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2603:26  */
  assign n8264_o = 1'b0 ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2611:38  */
  assign n8267_o = csr[433];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2617:46  */
  assign n8273_o = csr[432];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2617:40  */
  assign n8275_o = {3'b000, n8273_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2623:38  */
  assign n8283_o = 1'b0 ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2624:38  */
  assign n8285_o = csr[431];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:395:5  */
  always @(posedge clk_i or posedge n2790_o)
    if (n2790_o)
      n8288_q <= 1'b0;
    else
      n8288_q <= n2877_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:395:5  */
  always @(posedge clk_i or posedge n2790_o)
    if (n2790_o)
      n8289_q <= n2883_o;
    else
      n8289_q <= n2878_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:388:5  */
  assign n8290_o = {n8288_q, n2903_o, n2907_o, n3824_o, n8289_q};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:388:5  */
  assign n8291_o = {prefetch_buffer_n2_prefetch_buffer_inst_n2964, prefetch_buffer_n1_prefetch_buffer_inst_n2949, n3094_o, n3086_o, prefetch_buffer_n1_prefetch_buffer_inst_n2948, prefetch_buffer_n2_prefetch_buffer_inst_n2963, prefetch_buffer_n2_prefetch_buffer_inst_n2961, prefetch_buffer_n1_prefetch_buffer_inst_n2946, n2940_o, n2932_o, n2914_o, n2920_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:520:7  */
  always @(posedge clk_i)
    n8292_q <= n2987_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:520:7  */
  assign n8293_o = {n3078_o, neorv32_cpu_decompressor_inst_true_neorv32_cpu_decompressor_inst_n3097, neorv32_cpu_decompressor_inst_true_neorv32_cpu_decompressor_inst_n3098, n3106_o, n3077_o, n3029_o, n8292_q};
  assign n8294_o = {n3456_o, n3451_o, 1'b0, 1'b0, 1'b0, n3446_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:671:5  */
  always @(posedge clk_i or posedge n3281_o)
    if (n3281_o)
      n8295_q <= 1'b1;
    else
      n8295_q <= n3297_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:671:5  */
  always @(posedge clk_i or posedge n3281_o)
    if (n3281_o)
      n8296_q <= n3362_o;
    else
      n8296_q <= n3343_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:671:5  */
  always @(posedge clk_i or posedge n3281_o)
    if (n3281_o)
      n8297_q <= 32'b00000000000000000000000000000000;
    else
      n8297_q <= n3341_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:671:5  */
  assign n8298_o = execute_engine[116:85];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:671:5  */
  assign n8299_o = n3308_o ? n3317_o : n8298_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:671:5  */
  always @(posedge clk_i or posedge n3281_o)
    if (n3281_o)
      n8300_q <= 32'b11111111111111110000000000000000;
    else
      n8300_q <= n8299_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:671:5  */
  always @(posedge clk_i or posedge n3281_o)
    if (n3281_o)
      n8301_q <= 1'b0;
    else
      n8301_q <= n3300_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:671:5  */
  always @(posedge clk_i or posedge n3281_o)
    if (n3281_o)
      n8302_q <= 1'b0;
    else
      n8302_q <= n3299_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:671:5  */
  always @(posedge clk_i or posedge n3281_o)
    if (n3281_o)
      n8303_q <= n3361_o;
    else
      n8303_q <= n3342_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:671:5  */
  always @(posedge clk_i or posedge n3281_o)
    if (n3281_o)
      n8304_q <= 4'b0000;
    else
      n8304_q <= n3294_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:658:5  */
  assign n8305_o = {n3832_o, n8295_q, n3831_o, n8296_q, 28'b0000000000000000000000000000, n3380_o, n8297_q, n3830_o, n3829_o, n8300_q, n3278_o, n3828_o, n8301_q, n3827_o, n8302_q, n3826_o, n8303_q, n3825_o, n8304_q};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1602:5  */
  always @(posedge clk_i)
    n8306_q <= n5367_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1561:5  */
  always @(posedge clk_i or posedge n5128_o)
    if (n5128_o)
      n8307_q <= 1'b0;
    else
      n8307_q <= n5151_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1464:5  */
  always @(posedge clk_i or posedge n4842_o)
    if (n4842_o)
      n8308_q <= n5123_o;
    else
      n8308_q <= n5118_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1464:5  */
  always @(posedge clk_i or posedge n4842_o)
    if (n4842_o)
      n8309_q <= 11'b00000000000;
    else
      n8309_q <= n5117_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1460:5  */
  assign n8310_o = {n3838_o, n4839_o, n3836_o, n3834_o, n3833_o, n8307_q, n5263_o, n8306_q, n5253_o, n8308_q, n5188_o, n8309_q};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1460:5  */
  assign n8311_o = {n3866_o, n3857_o, n3855_o, n3853_o, n3864_o, n3851_o, n3849_o, n3861_o, n3488_o, n3847_o, n3845_o, n3843_o, n3842_o, n3841_o, n3858_o, n3840_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:671:5  */
  always @(posedge clk_i or posedge n3281_o)
    if (n3281_o)
      n8312_q <= 70'b0000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n8312_q <= ctrl_nxt;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2123:5  */
  always @(posedge clk_i)
    n8313_q <= n6716_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2123:5  */
  always @(posedge clk_i)
    n8314_q <= n5705_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1706:5  */
  always @(posedge clk_i or posedge n5393_o)
    if (n5393_o)
      n8315_q <= 32'b00000000000000000000000000000000;
    else
      n8315_q <= 32'b00000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1706:5  */
  always @(posedge clk_i or posedge n5393_o)
    if (n5393_o)
      n8316_q <= n5641_o;
    else
      n8316_q <= n5628_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1706:5  */
  always @(posedge clk_i or posedge n5393_o)
    if (n5393_o)
      n8317_q <= n5640_o;
    else
      n8317_q <= n5627_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1706:5  */
  always @(posedge clk_i or posedge n5393_o)
    if (n5393_o)
      n8318_q <= n5639_o;
    else
      n8318_q <= n5626_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1706:5  */
  always @(posedge clk_i or posedge n5393_o)
    if (n5393_o)
      n8319_q <= 1'b0;
    else
      n8319_q <= n5430_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:1673:5  */
  assign n8320_o = {n8315_q, 4'b0010, n8267_o, 6'b000000, 1'b0, 1'b0, 1'b1, 2'b00, n8275_o, 1'b0, 4'b0000, 1'b1, 1'b0, 1'b0, n8283_o, n8285_o, 1'b0, 1'b0, n8316_q, 4'b0100, 12'b000000000000, n8244_o, 1'b0, 1'b0, n8249_o, 1'b0, 1'b1, 1'b0, n8254_o, 1'b0, 1'b1, 1'b0, n8258_o, n8261_o, n8317_q, n5650_o, n8318_q, n8313_q, n5390_o, n3868_o, n8314_q, n3867_o, n8319_q, n3458_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2488:5  */
  always @(posedge clk_i)
    n8322_q <= n8082_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n8000_o)
    if (n8000_o)
      n8323_q <= 1'b0;
    else
      n8323_q <= n8009_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n8000_o)
    if (n8000_o)
      n8324_q <= 32'b00000000000000000000000000000000;
    else
      n8324_q <= n8016_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n8000_o)
    if (n8000_o)
      n8325_q <= 32'b00000000000000000000000000000000;
    else
      n8325_q <= n8008_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7960_o)
    if (n7960_o)
      n8326_q <= 1'b0;
    else
      n8326_q <= n7969_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7960_o)
    if (n7960_o)
      n8327_q <= 32'b00000000000000000000000000000000;
    else
      n8327_q <= n7976_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7960_o)
    if (n7960_o)
      n8328_q <= 32'b00000000000000000000000000000000;
    else
      n8328_q <= n7968_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7920_o)
    if (n7920_o)
      n8329_q <= 1'b0;
    else
      n8329_q <= n7929_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7920_o)
    if (n7920_o)
      n8330_q <= 32'b00000000000000000000000000000000;
    else
      n8330_q <= n7936_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7920_o)
    if (n7920_o)
      n8331_q <= 32'b00000000000000000000000000000000;
    else
      n8331_q <= n7928_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7880_o)
    if (n7880_o)
      n8332_q <= 1'b0;
    else
      n8332_q <= n7889_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7880_o)
    if (n7880_o)
      n8333_q <= 32'b00000000000000000000000000000000;
    else
      n8333_q <= n7896_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7880_o)
    if (n7880_o)
      n8334_q <= 32'b00000000000000000000000000000000;
    else
      n8334_q <= n7888_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7840_o)
    if (n7840_o)
      n8335_q <= 1'b0;
    else
      n8335_q <= n7849_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7840_o)
    if (n7840_o)
      n8336_q <= 32'b00000000000000000000000000000000;
    else
      n8336_q <= n7856_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7840_o)
    if (n7840_o)
      n8337_q <= 32'b00000000000000000000000000000000;
    else
      n8337_q <= n7848_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7800_o)
    if (n7800_o)
      n8338_q <= 1'b0;
    else
      n8338_q <= n7809_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7800_o)
    if (n7800_o)
      n8339_q <= 32'b00000000000000000000000000000000;
    else
      n8339_q <= n7816_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7800_o)
    if (n7800_o)
      n8340_q <= 32'b00000000000000000000000000000000;
    else
      n8340_q <= n7808_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7760_o)
    if (n7760_o)
      n8341_q <= 1'b0;
    else
      n8341_q <= n7769_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7760_o)
    if (n7760_o)
      n8342_q <= 32'b00000000000000000000000000000000;
    else
      n8342_q <= n7776_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7760_o)
    if (n7760_o)
      n8343_q <= 32'b00000000000000000000000000000000;
    else
      n8343_q <= n7768_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7720_o)
    if (n7720_o)
      n8344_q <= 1'b0;
    else
      n8344_q <= n7729_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7720_o)
    if (n7720_o)
      n8345_q <= 32'b00000000000000000000000000000000;
    else
      n8345_q <= n7736_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7720_o)
    if (n7720_o)
      n8346_q <= 32'b00000000000000000000000000000000;
    else
      n8346_q <= n7728_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7680_o)
    if (n7680_o)
      n8347_q <= 1'b0;
    else
      n8347_q <= n7689_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7680_o)
    if (n7680_o)
      n8348_q <= 32'b00000000000000000000000000000000;
    else
      n8348_q <= n7696_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7680_o)
    if (n7680_o)
      n8349_q <= 32'b00000000000000000000000000000000;
    else
      n8349_q <= n7688_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7640_o)
    if (n7640_o)
      n8350_q <= 1'b0;
    else
      n8350_q <= n7649_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7640_o)
    if (n7640_o)
      n8351_q <= 32'b00000000000000000000000000000000;
    else
      n8351_q <= n7656_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7640_o)
    if (n7640_o)
      n8352_q <= 32'b00000000000000000000000000000000;
    else
      n8352_q <= n7648_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7600_o)
    if (n7600_o)
      n8353_q <= 1'b0;
    else
      n8353_q <= n7609_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7600_o)
    if (n7600_o)
      n8354_q <= 32'b00000000000000000000000000000000;
    else
      n8354_q <= n7616_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7600_o)
    if (n7600_o)
      n8355_q <= 32'b00000000000000000000000000000000;
    else
      n8355_q <= n7608_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7560_o)
    if (n7560_o)
      n8356_q <= 1'b0;
    else
      n8356_q <= n7569_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7560_o)
    if (n7560_o)
      n8357_q <= 32'b00000000000000000000000000000000;
    else
      n8357_q <= n7576_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7560_o)
    if (n7560_o)
      n8358_q <= 32'b00000000000000000000000000000000;
    else
      n8358_q <= n7568_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7520_o)
    if (n7520_o)
      n8359_q <= 1'b0;
    else
      n8359_q <= n7529_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7520_o)
    if (n7520_o)
      n8360_q <= 32'b00000000000000000000000000000000;
    else
      n8360_q <= n7536_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7520_o)
    if (n7520_o)
      n8361_q <= 32'b00000000000000000000000000000000;
    else
      n8361_q <= n7528_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7480_o)
    if (n7480_o)
      n8362_q <= 1'b0;
    else
      n8362_q <= n7489_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7480_o)
    if (n7480_o)
      n8363_q <= 32'b00000000000000000000000000000000;
    else
      n8363_q <= n7496_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7480_o)
    if (n7480_o)
      n8364_q <= 32'b00000000000000000000000000000000;
    else
      n8364_q <= n7488_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7440_o)
    if (n7440_o)
      n8365_q <= 1'b0;
    else
      n8365_q <= n7449_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7440_o)
    if (n7440_o)
      n8366_q <= 32'b00000000000000000000000000000000;
    else
      n8366_q <= n7456_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7440_o)
    if (n7440_o)
      n8367_q <= 32'b00000000000000000000000000000000;
    else
      n8367_q <= n7448_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7400_o)
    if (n7400_o)
      n8368_q <= 1'b0;
    else
      n8368_q <= n7409_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7400_o)
    if (n7400_o)
      n8369_q <= 32'b00000000000000000000000000000000;
    else
      n8369_q <= n7416_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7400_o)
    if (n7400_o)
      n8370_q <= 32'b00000000000000000000000000000000;
    else
      n8370_q <= n7408_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7360_o)
    if (n7360_o)
      n8371_q <= 1'b0;
    else
      n8371_q <= n7369_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7360_o)
    if (n7360_o)
      n8372_q <= 32'b00000000000000000000000000000000;
    else
      n8372_q <= n7376_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7360_o)
    if (n7360_o)
      n8373_q <= 32'b00000000000000000000000000000000;
    else
      n8373_q <= n7368_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7320_o)
    if (n7320_o)
      n8374_q <= 1'b0;
    else
      n8374_q <= n7329_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7320_o)
    if (n7320_o)
      n8375_q <= 32'b00000000000000000000000000000000;
    else
      n8375_q <= n7336_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7320_o)
    if (n7320_o)
      n8376_q <= 32'b00000000000000000000000000000000;
    else
      n8376_q <= n7328_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7280_o)
    if (n7280_o)
      n8377_q <= 1'b0;
    else
      n8377_q <= n7289_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7280_o)
    if (n7280_o)
      n8378_q <= 32'b00000000000000000000000000000000;
    else
      n8378_q <= n7296_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7280_o)
    if (n7280_o)
      n8379_q <= 32'b00000000000000000000000000000000;
    else
      n8379_q <= n7288_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7240_o)
    if (n7240_o)
      n8380_q <= 1'b0;
    else
      n8380_q <= n7249_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7240_o)
    if (n7240_o)
      n8381_q <= 32'b00000000000000000000000000000000;
    else
      n8381_q <= n7256_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7240_o)
    if (n7240_o)
      n8382_q <= 32'b00000000000000000000000000000000;
    else
      n8382_q <= n7248_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7200_o)
    if (n7200_o)
      n8383_q <= 1'b0;
    else
      n8383_q <= n7209_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7200_o)
    if (n7200_o)
      n8384_q <= 32'b00000000000000000000000000000000;
    else
      n8384_q <= n7216_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7200_o)
    if (n7200_o)
      n8385_q <= 32'b00000000000000000000000000000000;
    else
      n8385_q <= n7208_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7160_o)
    if (n7160_o)
      n8386_q <= 1'b0;
    else
      n8386_q <= n7169_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7160_o)
    if (n7160_o)
      n8387_q <= 32'b00000000000000000000000000000000;
    else
      n8387_q <= n7176_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7160_o)
    if (n7160_o)
      n8388_q <= 32'b00000000000000000000000000000000;
    else
      n8388_q <= n7168_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7120_o)
    if (n7120_o)
      n8389_q <= 1'b0;
    else
      n8389_q <= n7129_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7120_o)
    if (n7120_o)
      n8390_q <= 32'b00000000000000000000000000000000;
    else
      n8390_q <= n7136_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7120_o)
    if (n7120_o)
      n8391_q <= 32'b00000000000000000000000000000000;
    else
      n8391_q <= n7128_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7080_o)
    if (n7080_o)
      n8392_q <= 1'b0;
    else
      n8392_q <= n7089_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7080_o)
    if (n7080_o)
      n8393_q <= 32'b00000000000000000000000000000000;
    else
      n8393_q <= n7096_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7080_o)
    if (n7080_o)
      n8394_q <= 32'b00000000000000000000000000000000;
    else
      n8394_q <= n7088_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7040_o)
    if (n7040_o)
      n8395_q <= 1'b0;
    else
      n8395_q <= n7049_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7040_o)
    if (n7040_o)
      n8396_q <= 32'b00000000000000000000000000000000;
    else
      n8396_q <= n7056_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7040_o)
    if (n7040_o)
      n8397_q <= 32'b00000000000000000000000000000000;
    else
      n8397_q <= n7048_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7000_o)
    if (n7000_o)
      n8398_q <= 1'b0;
    else
      n8398_q <= n7009_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7000_o)
    if (n7000_o)
      n8399_q <= 32'b00000000000000000000000000000000;
    else
      n8399_q <= n7016_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n7000_o)
    if (n7000_o)
      n8400_q <= 32'b00000000000000000000000000000000;
    else
      n8400_q <= n7008_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6960_o)
    if (n6960_o)
      n8401_q <= 1'b0;
    else
      n8401_q <= n6969_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6960_o)
    if (n6960_o)
      n8402_q <= 32'b00000000000000000000000000000000;
    else
      n8402_q <= n6976_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6960_o)
    if (n6960_o)
      n8403_q <= 32'b00000000000000000000000000000000;
    else
      n8403_q <= n6968_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6920_o)
    if (n6920_o)
      n8404_q <= 1'b0;
    else
      n8404_q <= n6929_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6920_o)
    if (n6920_o)
      n8405_q <= 32'b00000000000000000000000000000000;
    else
      n8405_q <= n6936_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6920_o)
    if (n6920_o)
      n8406_q <= 32'b00000000000000000000000000000000;
    else
      n8406_q <= n6928_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6880_o)
    if (n6880_o)
      n8407_q <= 1'b0;
    else
      n8407_q <= n6889_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6880_o)
    if (n6880_o)
      n8408_q <= 32'b00000000000000000000000000000000;
    else
      n8408_q <= n6896_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6880_o)
    if (n6880_o)
      n8409_q <= 32'b00000000000000000000000000000000;
    else
      n8409_q <= n6888_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6840_o)
    if (n6840_o)
      n8410_q <= 1'b0;
    else
      n8410_q <= n6849_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6840_o)
    if (n6840_o)
      n8411_q <= 32'b00000000000000000000000000000000;
    else
      n8411_q <= n6856_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6840_o)
    if (n6840_o)
      n8412_q <= 32'b00000000000000000000000000000000;
    else
      n8412_q <= n6848_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6800_o)
    if (n6800_o)
      n8413_q <= 1'b0;
    else
      n8413_q <= n6809_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6800_o)
    if (n6800_o)
      n8414_q <= 32'b00000000000000000000000000000000;
    else
      n8414_q <= n6816_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6800_o)
    if (n6800_o)
      n8415_q <= 32'b00000000000000000000000000000000;
    else
      n8415_q <= n6808_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6760_o)
    if (n6760_o)
      n8416_q <= 1'b0;
    else
      n8416_q <= n6769_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6760_o)
    if (n6760_o)
      n8417_q <= 32'b00000000000000000000000000000000;
    else
      n8417_q <= n6776_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2433:7  */
  always @(posedge clk_i or posedge n6760_o)
    if (n6760_o)
      n8418_q <= 32'b00000000000000000000000000000000;
    else
      n8418_q <= n6768_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:7  */
  assign n8419_o = {n8416_q, n8413_q, n8410_q, n8407_q, n8404_q, n8401_q, n8398_q, n8395_q, n8392_q, n8389_q, n8386_q, n8383_q, n8380_q, n8377_q, n8374_q, n8371_q, n8368_q, n8365_q, n8362_q, n8359_q, n8356_q, n8353_q, n8350_q, n8347_q, n8344_q, n8341_q, n8338_q, n8335_q, n8332_q, n8329_q, n8326_q, n8323_q, n6793_o, n6833_o, n6873_o, n6913_o, n6953_o, n6993_o, n7033_o, n7073_o, n7113_o, n7153_o, n7193_o, n7233_o, n7273_o, n7313_o, n7353_o, n7393_o, n7433_o, n7473_o, n7513_o, n7553_o, n7593_o, n7633_o, n7673_o, n7713_o, n7753_o, n7793_o, n7833_o, n7873_o, n7913_o, n7953_o, n7993_o, n8033_o, n8417_q, n8414_q, n8411_q, n8408_q, n8405_q, n8402_q, n8399_q, n8396_q, n8393_q, n8390_q, n8387_q, n8384_q, n8381_q, n8378_q, n8375_q, n8372_q, n8369_q, n8366_q, n8363_q, n8360_q, n8357_q, n8354_q, n8351_q, n8348_q, n8345_q, n8342_q, n8339_q, n8336_q, n8333_q, n8330_q, n8327_q, n8324_q, n8418_q, n8415_q, n8412_q, n8409_q, n8406_q, n8403_q, n8400_q, n8397_q, n8394_q, n8391_q, n8388_q, n8385_q, n8382_q, n8379_q, n8376_q, n8373_q, n8370_q, n8367_q, n8364_q, n8361_q, n8358_q, n8355_q, n8352_q, n8349_q, n8346_q, n8343_q, n8340_q, n8337_q, n8334_q, n8331_q, n8328_q, n8325_q, n8322_q, n6757_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:7  */
  assign n8420_o = {n8040_o, n8046_o, n8050_o, n8051_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:7  */
  assign n8421_o = {n8043_o, n8048_o, n8052_o, n8053_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2429:7  */
  assign n8422_o = {n8195_o, n8187_o, n8183_o, n8170_o, n8161_o, n8153_o, n8143_o, n8137_o, n8130_o, n8124_o, n8114_o, n8104_o, n8096_o, 1'b0, n8089_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2536:5  */
  always @(posedge clk_i or posedge n8198_o)
    if (n8198_o)
      n8423_q <= 1'b0;
    else
      n8423_q <= 1'b0;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2536:5  */
  always @(posedge clk_i or posedge n8198_o)
    if (n8198_o)
      n8424_q <= 2'b00;
    else
      n8424_q <= 2'b00;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2533:5  */
  assign n8425_o = {n8423_q, n3869_o, n8241_o, n8237_o, n8233_o, n8221_o, n8213_o, n8424_q};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2533:5  */
  assign n8426_o = {n3419_o, n3418_o, n3417_o, n3416_o, n3415_o, n3414_o, n3413_o, n3412_o, n3408_o, n3407_o, n3406_o, n3405_o, n3404_o, n3403_o, n3402_o, n3401_o, n3400_o, n3399_o, n3398_o, n3397_o, n3396_o, n3395_o, n3394_o, n3393_o, n3392_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:609:5  */
  always @(posedge clk_i)
    n8427_q <= n3263_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8428_o = n6743_o[4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8429_o = ~n8428_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8430_o = n6743_o[3];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8431_o = ~n8430_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8432_o = n8429_o & n8431_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8433_o = n8429_o & n8430_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8434_o = n8428_o & n8431_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8435_o = n8428_o & n8430_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8436_o = n6743_o[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8437_o = ~n8436_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8438_o = n8432_o & n8437_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8439_o = n8432_o & n8436_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8440_o = n8433_o & n8437_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8441_o = n8433_o & n8436_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8442_o = n8434_o & n8437_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8443_o = n8434_o & n8436_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8444_o = n8435_o & n8437_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8445_o = n8435_o & n8436_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8446_o = n6743_o[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8447_o = ~n8446_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8448_o = n8438_o & n8447_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8449_o = n8438_o & n8446_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8450_o = n8439_o & n8447_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8451_o = n8439_o & n8446_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8452_o = n8440_o & n8447_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8453_o = n8440_o & n8446_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8454_o = n8441_o & n8447_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8455_o = n8441_o & n8446_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8456_o = n8442_o & n8447_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8457_o = n8442_o & n8446_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8458_o = n8443_o & n8447_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8459_o = n8443_o & n8446_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8460_o = n8444_o & n8447_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8461_o = n8444_o & n8446_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8462_o = n8445_o & n8447_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8463_o = n8445_o & n8446_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8464_o = n6743_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8465_o = ~n8464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8466_o = n8448_o & n8465_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8467_o = n8448_o & n8464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8468_o = n8449_o & n8465_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8469_o = n8449_o & n8464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8470_o = n8450_o & n8465_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8471_o = n8450_o & n8464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8472_o = n8451_o & n8465_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8473_o = n8451_o & n8464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8474_o = n8452_o & n8465_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8475_o = n8452_o & n8464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8476_o = n8453_o & n8465_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8477_o = n8453_o & n8464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8478_o = n8454_o & n8465_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8479_o = n8454_o & n8464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8480_o = n8455_o & n8465_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8481_o = n8455_o & n8464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8482_o = n8456_o & n8465_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8483_o = n8456_o & n8464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8484_o = n8457_o & n8465_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8485_o = n8457_o & n8464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8486_o = n8458_o & n8465_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8487_o = n8458_o & n8464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8488_o = n8459_o & n8465_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8489_o = n8459_o & n8464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8490_o = n8460_o & n8465_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8491_o = n8460_o & n8464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8492_o = n8461_o & n8465_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8493_o = n8461_o & n8464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8494_o = n8462_o & n8465_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8495_o = n8462_o & n8464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8496_o = n8463_o & n8465_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8497_o = n8463_o & n8464_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2427:5  */
  assign n8498_o = n6734_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8499_o = n8466_o ? 1'b1 : n8498_o;
  assign n8500_o = n6734_o[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8501_o = n8467_o ? 1'b1 : n8500_o;
  assign n8502_o = n6734_o[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8503_o = n8468_o ? 1'b1 : n8502_o;
  assign n8504_o = n6734_o[3];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8505_o = n8469_o ? 1'b1 : n8504_o;
  assign n8506_o = n6734_o[4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8507_o = n8470_o ? 1'b1 : n8506_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2427:5  */
  assign n8508_o = n6734_o[5];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8509_o = n8471_o ? 1'b1 : n8508_o;
  assign n8510_o = n6734_o[6];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8511_o = n8472_o ? 1'b1 : n8510_o;
  assign n8512_o = n6734_o[7];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8513_o = n8473_o ? 1'b1 : n8512_o;
  assign n8514_o = n6734_o[8];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8515_o = n8474_o ? 1'b1 : n8514_o;
  assign n8516_o = n6734_o[9];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8517_o = n8475_o ? 1'b1 : n8516_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2427:5  */
  assign n8518_o = n6734_o[10];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8519_o = n8476_o ? 1'b1 : n8518_o;
  assign n8520_o = n6734_o[11];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8521_o = n8477_o ? 1'b1 : n8520_o;
  assign n8522_o = n6734_o[12];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8523_o = n8478_o ? 1'b1 : n8522_o;
  assign n8524_o = n6734_o[13];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8525_o = n8479_o ? 1'b1 : n8524_o;
  assign n8526_o = n6734_o[14];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8527_o = n8480_o ? 1'b1 : n8526_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2427:5  */
  assign n8528_o = n6734_o[15];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8529_o = n8481_o ? 1'b1 : n8528_o;
  assign n8530_o = n6734_o[16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8531_o = n8482_o ? 1'b1 : n8530_o;
  assign n8532_o = n6734_o[17];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8533_o = n8483_o ? 1'b1 : n8532_o;
  assign n8534_o = n6734_o[18];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8535_o = n8484_o ? 1'b1 : n8534_o;
  assign n8536_o = n6734_o[19];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8537_o = n8485_o ? 1'b1 : n8536_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2427:5  */
  assign n8538_o = n6734_o[20];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8539_o = n8486_o ? 1'b1 : n8538_o;
  assign n8540_o = n6734_o[21];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8541_o = n8487_o ? 1'b1 : n8540_o;
  assign n8542_o = n6734_o[22];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8543_o = n8488_o ? 1'b1 : n8542_o;
  assign n8544_o = n6734_o[23];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8545_o = n8489_o ? 1'b1 : n8544_o;
  assign n8546_o = n6734_o[24];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8547_o = n8490_o ? 1'b1 : n8546_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2427:5  */
  assign n8548_o = n6734_o[25];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8549_o = n8491_o ? 1'b1 : n8548_o;
  assign n8550_o = n6734_o[26];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8551_o = n8492_o ? 1'b1 : n8550_o;
  assign n8552_o = n6734_o[27];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8553_o = n8493_o ? 1'b1 : n8552_o;
  assign n8554_o = n6734_o[28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8555_o = n8494_o ? 1'b1 : n8554_o;
  assign n8556_o = n6734_o[29];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8557_o = n8495_o ? 1'b1 : n8556_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2427:5  */
  assign n8558_o = n6734_o[30];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8559_o = n8496_o ? 1'b1 : n8558_o;
  assign n8560_o = n6734_o[31];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:9  */
  assign n8561_o = n8497_o ? 1'b1 : n8560_o;
  assign n8562_o = {n8561_o, n8559_o, n8557_o, n8555_o, n8553_o, n8551_o, n8549_o, n8547_o, n8545_o, n8543_o, n8541_o, n8539_o, n8537_o, n8535_o, n8533_o, n8531_o, n8529_o, n8527_o, n8525_o, n8523_o, n8521_o, n8519_o, n8517_o, n8515_o, n8513_o, n8511_o, n8509_o, n8507_o, n8505_o, n8503_o, n8501_o, n8499_o};
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8563_o = n6748_o[4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8564_o = ~n8563_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8565_o = n6748_o[3];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8566_o = ~n8565_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8567_o = n8564_o & n8566_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8568_o = n8564_o & n8565_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8569_o = n8563_o & n8566_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8570_o = n8563_o & n8565_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8571_o = n6748_o[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8572_o = ~n8571_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8573_o = n8567_o & n8572_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8574_o = n8567_o & n8571_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8575_o = n8568_o & n8572_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8576_o = n8568_o & n8571_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8577_o = n8569_o & n8572_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8578_o = n8569_o & n8571_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8579_o = n8570_o & n8572_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8580_o = n8570_o & n8571_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8581_o = n6748_o[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8582_o = ~n8581_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8583_o = n8573_o & n8582_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8584_o = n8573_o & n8581_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8585_o = n8574_o & n8582_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8586_o = n8574_o & n8581_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8587_o = n8575_o & n8582_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8588_o = n8575_o & n8581_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8589_o = n8576_o & n8582_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8590_o = n8576_o & n8581_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8591_o = n8577_o & n8582_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8592_o = n8577_o & n8581_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8593_o = n8578_o & n8582_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8594_o = n8578_o & n8581_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8595_o = n8579_o & n8582_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8596_o = n8579_o & n8581_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8597_o = n8580_o & n8582_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8598_o = n8580_o & n8581_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8599_o = n6748_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8600_o = ~n8599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8601_o = n8583_o & n8600_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8602_o = n8583_o & n8599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8603_o = n8584_o & n8600_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8604_o = n8584_o & n8599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8605_o = n8585_o & n8600_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8606_o = n8585_o & n8599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8607_o = n8586_o & n8600_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8608_o = n8586_o & n8599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8609_o = n8587_o & n8600_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8610_o = n8587_o & n8599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8611_o = n8588_o & n8600_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8612_o = n8588_o & n8599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8613_o = n8589_o & n8600_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8614_o = n8589_o & n8599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8615_o = n8590_o & n8600_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8616_o = n8590_o & n8599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8617_o = n8591_o & n8600_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8618_o = n8591_o & n8599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8619_o = n8592_o & n8600_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8620_o = n8592_o & n8599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8621_o = n8593_o & n8600_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8622_o = n8593_o & n8599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8623_o = n8594_o & n8600_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8624_o = n8594_o & n8599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8625_o = n8595_o & n8600_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8626_o = n8595_o & n8599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8627_o = n8596_o & n8600_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8628_o = n8596_o & n8599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8629_o = n8597_o & n8600_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8630_o = n8597_o & n8599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8631_o = n8598_o & n8600_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8632_o = n8598_o & n8599_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2416:19  */
  assign n8633_o = n6735_o[0];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8634_o = n8601_o ? 1'b1 : n8633_o;
  assign n8635_o = n6735_o[1];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8636_o = n8602_o ? 1'b1 : n8635_o;
  assign n8637_o = n6735_o[2];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8638_o = n8603_o ? 1'b1 : n8637_o;
  assign n8639_o = n6735_o[3];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8640_o = n8604_o ? 1'b1 : n8639_o;
  assign n8641_o = n6735_o[4];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8642_o = n8605_o ? 1'b1 : n8641_o;
  assign n8643_o = n6735_o[5];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8644_o = n8606_o ? 1'b1 : n8643_o;
  assign n8645_o = n6735_o[6];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8646_o = n8607_o ? 1'b1 : n8645_o;
  assign n8647_o = n6735_o[7];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8648_o = n8608_o ? 1'b1 : n8647_o;
  assign n8649_o = n6735_o[8];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8650_o = n8609_o ? 1'b1 : n8649_o;
  assign n8651_o = n6735_o[9];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8652_o = n8610_o ? 1'b1 : n8651_o;
  assign n8653_o = n6735_o[10];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8654_o = n8611_o ? 1'b1 : n8653_o;
  assign n8655_o = n6735_o[11];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8656_o = n8612_o ? 1'b1 : n8655_o;
  assign n8657_o = n6735_o[12];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8658_o = n8613_o ? 1'b1 : n8657_o;
  assign n8659_o = n6735_o[13];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8660_o = n8614_o ? 1'b1 : n8659_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2121:3  */
  assign n8661_o = n6735_o[14];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8662_o = n8615_o ? 1'b1 : n8661_o;
  assign n8663_o = n6735_o[15];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8664_o = n8616_o ? 1'b1 : n8663_o;
  assign n8665_o = n6735_o[16];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8666_o = n8617_o ? 1'b1 : n8665_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2088:5  */
  assign n8667_o = n6735_o[17];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8668_o = n8618_o ? 1'b1 : n8667_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2089:7  */
  assign n8669_o = n6735_o[18];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8670_o = n8619_o ? 1'b1 : n8669_o;
  assign n8671_o = n6735_o[19];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8672_o = n8620_o ? 1'b1 : n8671_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2089:19  */
  assign n8673_o = n6735_o[20];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8674_o = n8621_o ? 1'b1 : n8673_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2088:50  */
  assign n8675_o = n6735_o[21];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8676_o = n8622_o ? 1'b1 : n8675_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2088:31  */
  assign n8677_o = n6735_o[22];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8678_o = n8623_o ? 1'b1 : n8677_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2088:17  */
  assign n8679_o = n6735_o[23];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8680_o = n8624_o ? 1'b1 : n8679_o;
  assign n8681_o = n6735_o[24];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8682_o = n8625_o ? 1'b1 : n8681_o;
  assign n8683_o = n6735_o[25];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8684_o = n8626_o ? 1'b1 : n8683_o;
  assign n8685_o = n6735_o[26];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8686_o = n8627_o ? 1'b1 : n8685_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2016:7  */
  assign n8687_o = n6735_o[27];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8688_o = n8628_o ? 1'b1 : n8687_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2016:19  */
  assign n8689_o = n6735_o[28];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8690_o = n8629_o ? 1'b1 : n8689_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2016:47  */
  assign n8691_o = n6735_o[29];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8692_o = n8630_o ? 1'b1 : n8691_o;
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2015:63  */
  assign n8693_o = n6735_o[30];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8694_o = n8631_o ? 1'b1 : n8693_o;
  assign n8695_o = n6735_o[31];
  /* ../neorv32/rtl/core/neorv32_cpu_control.vhd:2418:9  */
  assign n8696_o = n8632_o ? 1'b1 : n8695_o;
  assign n8697_o = {n8696_o, n8694_o, n8692_o, n8690_o, n8688_o, n8686_o, n8684_o, n8682_o, n8680_o, n8678_o, n8676_o, n8674_o, n8672_o, n8670_o, n8668_o, n8666_o, n8664_o, n8662_o, n8660_o, n8658_o, n8656_o, n8654_o, n8652_o, n8650_o, n8648_o, n8646_o, n8644_o, n8642_o, n8640_o, n8638_o, n8636_o, n8634_o};
endmodule

module neorv32_sysinfo_5000000_0_1024_2048_4_64_1_4_64_0_0_0_c00c06f0c8f7e7aa711090f9c2d219a9079d700c
  (input  clk_i,
   input  [31:0] addr_i,
   input  rden_i,
   input  wren_i,
   output [31:0] data_o,
   output ack_o,
   output err_o);
  wire acc_en;
  wire rden;
  wire wren;
  wire [2:0] addr;
  wire [255:0] sysinfo;
  wire [3:0] n2619_o;
  wire n2621_o;
  wire n2622_o;
  wire n2624_o;
  wire n2625_o;
  wire [2:0] n2627_o;
  wire [3:0] n2685_o;
  wire [3:0] n2690_o;
  wire [3:0] n2695_o;
  wire [3:0] n2699_o;
  wire [3:0] n2704_o;
  wire [3:0] n2709_o;
  wire [31:0] n2717_o;
  wire [31:0] n2721_o;
  wire [2:0] n2727_o;
  wire [31:0] n2731_o;
  wire [255:0] n2737_o;
  reg [31:0] n2738_q;
  reg n2739_q;
  reg n2740_q;
  wire [31:0] n2741_o;
  wire [31:0] n2742_o;
  wire [31:0] n2743_o;
  wire [31:0] n2744_o;
  wire [31:0] n2745_o;
  wire [31:0] n2746_o;
  wire [31:0] n2747_o;
  wire [31:0] n2748_o;
  wire [1:0] n2749_o;
  reg [31:0] n2750_o;
  wire [1:0] n2751_o;
  reg [31:0] n2752_o;
  wire n2753_o;
  wire [31:0] n2754_o;
  assign data_o = n2738_q;
  assign ack_o = n2739_q;
  assign err_o = n2740_q;
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:110:10  */
  assign acc_en = n2622_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:111:10  */
  assign rden = n2624_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:112:10  */
  assign wren = n2625_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:113:10  */
  assign addr = n2627_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:117:10  */
  assign sysinfo = n2737_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:123:29  */
  assign n2619_o = addr_i[8:5];
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:123:56  */
  assign n2621_o = n2619_o == 4'b1111;
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:123:17  */
  assign n2622_o = n2621_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:124:20  */
  assign n2624_o = acc_en & rden_i;
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:125:20  */
  assign n2625_o = acc_en & wren_i;
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:126:19  */
  assign n2627_o = addr_i[4:2];
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:172:101  */
  assign n2685_o = 1'b0 ? 4'b0110 : 4'b0000;
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:173:101  */
  assign n2690_o = 1'b0 ? 4'b0010 : 4'b0000;
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:174:101  */
  assign n2695_o = 1'b0 ? 4'b0000 : 4'b0000;
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:175:38  */
  assign n2699_o = 1'b0 ? 4'b0001 : 4'b0000;
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:177:98  */
  assign n2704_o = 1'b0 ? 4'b0110 : 4'b0000;
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:178:98  */
  assign n2709_o = 1'b0 ? 4'b0010 : 4'b0000;
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:189:71  */
  assign n2717_o = 1'b1 ? 32'b00000000000000000000010000000000 : 32'b00000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:192:71  */
  assign n2721_o = 1'b1 ? 32'b00000000000000000000100000000000 : 32'b00000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:204:27  */
  assign n2727_o = 3'b111 - addr;
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:203:7  */
  assign n2731_o = rden ? n2754_o : 32'b00000000000000000000000000000000;
  assign n2737_o = {32'b00000000010011000100101101000000, 32'b00000000000000000000000000000000, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 6'b000000, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 4'b0000, 4'b0000, n2709_o, n2704_o, n2699_o, n2695_o, n2690_o, n2685_o, 32'b00000000000000000000000000000000, 32'b10000000000000000000000000000000, n2717_o, n2721_o};
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:199:5  */
  always @(posedge clk_i)
    n2738_q <= n2731_o;
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:199:5  */
  always @(posedge clk_i)
    n2739_q <= rden;
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:199:5  */
  always @(posedge clk_i)
    n2740_q <= wren;
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:99:5  */
  assign n2741_o = sysinfo[31:0];
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:98:5  */
  assign n2742_o = sysinfo[63:32];
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:97:5  */
  assign n2743_o = sysinfo[95:64];
  assign n2744_o = sysinfo[127:96];
  assign n2745_o = sysinfo[159:128];
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:204:27  */
  assign n2746_o = sysinfo[191:160];
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:197:3  */
  assign n2747_o = sysinfo[223:192];
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:199:5  */
  assign n2748_o = sysinfo[255:224];
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:204:26  */
  assign n2749_o = n2727_o[1:0];
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:204:26  */
  always @*
    case (n2749_o)
      2'b00: n2750_o = n2741_o;
      2'b01: n2750_o = n2742_o;
      2'b10: n2750_o = n2743_o;
      2'b11: n2750_o = n2744_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:204:26  */
  assign n2751_o = n2727_o[1:0];
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:204:26  */
  always @*
    case (n2751_o)
      2'b00: n2752_o = n2745_o;
      2'b01: n2752_o = n2746_o;
      2'b10: n2752_o = n2747_o;
      2'b11: n2752_o = n2748_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:204:26  */
  assign n2753_o = n2727_o[2];
  /* ../neorv32/rtl/core/neorv32_sysinfo.vhd:204:26  */
  assign n2754_o = n2753_o ? n2752_o : n2750_o;
endmodule

module neorv32_uart_256_256_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  clk_i,
   input  rstn_i,
   input  [31:0] addr_i,
   input  rden_i,
   input  wren_i,
   input  [31:0] data_i,
   input  [7:0] clkgen_i,
   input  uart_rxd_i,
   input  uart_cts_i,
   output [31:0] data_o,
   output ack_o,
   output clkgen_en_o,
   output uart_txd_o,
   output uart_rts_o,
   output irq_rx_o,
   output irq_tx_o);
  wire acc_en;
  wire [31:0] addr;
  wire wren;
  wire rden;
  wire uart_clk;
  wire [20:0] ctrl;
  wire [29:0] tx_engine;
  wire [30:0] rx_engine;
  wire [21:0] rx_fifo;
  wire [21:0] tx_fifo;
  wire [5:0] n2106_o;
  wire n2108_o;
  wire n2109_o;
  wire n2111_o;
  wire [29:0] n2113_o;
  wire [31:0] n2115_o;
  wire n2116_o;
  wire n2117_o;
  wire n2119_o;
  wire n2132_o;
  wire n2133_o;
  wire n2134_o;
  wire n2135_o;
  wire [2:0] n2136_o;
  wire [9:0] n2137_o;
  wire n2138_o;
  wire n2139_o;
  wire n2140_o;
  wire n2141_o;
  wire n2142_o;
  wire [20:0] n2143_o;
  wire n2145_o;
  wire [20:0] n2147_o;
  wire n2152_o;
  wire n2154_o;
  wire n2155_o;
  wire n2156_o;
  wire n2157_o;
  wire [2:0] n2158_o;
  wire [9:0] n2159_o;
  wire n2160_o;
  wire n2161_o;
  wire n2162_o;
  wire n2163_o;
  wire n2164_o;
  wire n2165_o;
  wire n2166_o;
  wire n2167_o;
  wire n2168_o;
  wire n2169_o;
  wire n2170_o;
  wire n2171_o;
  wire n2172_o;
  wire n2173_o;
  wire n2174_o;
  wire n2175_o;
  wire n2176_o;
  wire n2177_o;
  wire n2178_o;
  wire [7:0] n2179_o;
  wire [26:0] n2180_o;
  wire [1:0] n2181_o;
  wire [7:0] n2182_o;
  wire [7:0] n2183_o;
  wire [18:0] n2184_o;
  wire [18:0] n2186_o;
  wire [1:0] n2188_o;
  wire [26:0] n2189_o;
  wire [26:0] n2191_o;
  wire [1:0] n2193_o;
  localparam [31:0] n2194_o = 32'b00000000000000000000000000000000;
  wire [2:0] n2196_o;
  wire [31:0] n2197_o;
  wire n2201_o;
  wire [2:0] n2202_o;
  wire n2206_o;
  wire tx_engine_fifo_inst_n2207;
  wire [7:0] n2208_o;
  wire n2209_o;
  wire tx_engine_fifo_inst_n2210;
  wire n2211_o;
  wire [7:0] tx_engine_fifo_inst_n2212;
  wire tx_engine_fifo_inst_n2213;
  wire tx_engine_fifo_inst_half_o;
  wire tx_engine_fifo_inst_free_o;
  wire [7:0] tx_engine_fifo_inst_rdata_o;
  wire tx_engine_fifo_inst_avail_o;
  wire n2223_o;
  wire n2224_o;
  wire n2225_o;
  wire n2226_o;
  wire n2227_o;
  wire [7:0] n2229_o;
  wire n2232_o;
  wire n2233_o;
  wire n2234_o;
  wire [2:0] n2237_o;
  wire n2239_o;
  wire n2240_o;
  wire n2244_o;
  wire n2245_o;
  wire n2246_o;
  wire n2247_o;
  wire n2248_o;
  wire n2249_o;
  wire n2250_o;
  wire n2251_o;
  wire n2252_o;
  wire n2253_o;
  wire n2254_o;
  wire n2257_o;
  wire rx_engine_fifo_inst_n2258;
  wire [7:0] n2259_o;
  wire n2260_o;
  wire rx_engine_fifo_inst_n2261;
  wire n2262_o;
  wire [7:0] rx_engine_fifo_inst_n2263;
  wire rx_engine_fifo_inst_n2264;
  wire rx_engine_fifo_inst_half_o;
  wire rx_engine_fifo_inst_free_o;
  wire [7:0] rx_engine_fifo_inst_rdata_o;
  wire rx_engine_fifo_inst_avail_o;
  wire n2274_o;
  wire n2275_o;
  wire n2276_o;
  wire n2277_o;
  wire n2278_o;
  wire [7:0] n2280_o;
  wire n2281_o;
  wire n2284_o;
  wire n2285_o;
  wire n2286_o;
  wire n2290_o;
  wire n2291_o;
  wire n2292_o;
  wire n2293_o;
  wire n2294_o;
  wire n2295_o;
  wire n2296_o;
  wire n2297_o;
  wire n2298_o;
  wire n2299_o;
  wire n2300_o;
  wire n2301_o;
  wire n2302_o;
  wire n2303_o;
  wire n2308_o;
  wire [1:0] n2309_o;
  wire n2311_o;
  wire [2:0] n2312_o;
  wire [9:0] n2313_o;
  wire [7:0] n2315_o;
  wire [8:0] n2317_o;
  wire n2318_o;
  wire [1:0] n2320_o;
  wire [1:0] n2321_o;
  wire n2323_o;
  wire n2324_o;
  wire n2325_o;
  wire n2326_o;
  wire n2327_o;
  wire n2328_o;
  wire [1:0] n2330_o;
  wire [1:0] n2331_o;
  wire n2333_o;
  wire [9:0] n2335_o;
  wire n2341_o;
  wire n2343_o;
  wire n2345_o;
  wire n2346_o;
  wire n2347_o;
  wire n2348_o;
  wire n2349_o;
  wire n2350_o;
  wire n2351_o;
  wire n2352_o;
  wire n2353_o;
  wire n2354_o;
  wire n2355_o;
  wire n2356_o;
  wire n2357_o;
  wire n2358_o;
  wire n2359_o;
  wire n2360_o;
  wire n2361_o;
  wire n2362_o;
  wire n2363_o;
  wire [9:0] n2364_o;
  wire [3:0] n2365_o;
  wire [3:0] n2367_o;
  wire [7:0] n2368_o;
  wire [8:0] n2370_o;
  wire [9:0] n2371_o;
  wire [9:0] n2373_o;
  wire [22:0] n2374_o;
  wire [12:0] n2375_o;
  wire [12:0] n2376_o;
  wire [12:0] n2377_o;
  wire [9:0] n2378_o;
  wire [9:0] n2379_o;
  wire [22:0] n2380_o;
  wire [22:0] n2381_o;
  wire [22:0] n2382_o;
  wire [3:0] n2384_o;
  wire n2390_o;
  wire n2392_o;
  wire n2394_o;
  wire n2395_o;
  wire n2396_o;
  wire n2397_o;
  wire n2398_o;
  wire n2399_o;
  wire n2400_o;
  wire [1:0] n2403_o;
  wire [1:0] n2404_o;
  wire n2405_o;
  wire n2407_o;
  wire [2:0] n2409_o;
  reg [1:0] n2410_o;
  wire [8:0] n2411_o;
  wire [8:0] n2412_o;
  reg [8:0] n2413_o;
  wire [3:0] n2414_o;
  wire [3:0] n2415_o;
  reg [3:0] n2416_o;
  wire [9:0] n2417_o;
  wire [9:0] n2418_o;
  reg [9:0] n2419_o;
  reg n2420_o;
  wire [26:0] n2421_o;
  wire [1:0] n2428_o;
  wire n2430_o;
  wire n2431_o;
  wire n2433_o;
  wire [2:0] n2434_o;
  wire n2436_o;
  wire n2437_o;
  wire n2441_o;
  wire n2442_o;
  wire [1:0] n2443_o;
  wire [1:0] n2444_o;
  wire [1:0] n2445_o;
  wire n2447_o;
  wire [1:0] n2448_o;
  wire [8:0] n2449_o;
  wire [9:0] n2451_o;
  wire [1:0] n2453_o;
  wire n2455_o;
  wire n2457_o;
  wire n2458_o;
  wire n2460_o;
  wire [9:0] n2462_o;
  wire n2468_o;
  wire n2470_o;
  wire n2472_o;
  wire n2473_o;
  wire n2474_o;
  wire n2475_o;
  wire n2476_o;
  wire n2477_o;
  wire n2478_o;
  wire n2479_o;
  wire n2480_o;
  wire n2481_o;
  wire n2482_o;
  wire n2483_o;
  wire n2484_o;
  wire n2485_o;
  wire n2486_o;
  wire n2487_o;
  wire n2488_o;
  wire n2489_o;
  wire n2490_o;
  wire [9:0] n2491_o;
  wire [3:0] n2492_o;
  wire [3:0] n2494_o;
  wire n2495_o;
  wire [8:0] n2496_o;
  wire [9:0] n2497_o;
  wire [9:0] n2498_o;
  wire [9:0] n2500_o;
  wire [23:0] n2501_o;
  wire [13:0] n2502_o;
  wire [13:0] n2503_o;
  wire [13:0] n2504_o;
  wire [9:0] n2505_o;
  wire [9:0] n2506_o;
  wire [23:0] n2507_o;
  wire [23:0] n2508_o;
  wire [23:0] n2509_o;
  wire [3:0] n2511_o;
  wire n2517_o;
  wire n2519_o;
  wire n2521_o;
  wire n2522_o;
  wire n2523_o;
  wire n2524_o;
  wire n2525_o;
  wire n2526_o;
  wire n2527_o;
  wire n2530_o;
  wire n2531_o;
  wire n2532_o;
  wire n2534_o;
  wire [1:0] n2536_o;
  reg n2537_o;
  wire [9:0] n2538_o;
  wire [9:0] n2539_o;
  reg [9:0] n2540_o;
  wire [3:0] n2541_o;
  wire [3:0] n2542_o;
  reg [3:0] n2543_o;
  wire [9:0] n2544_o;
  wire [9:0] n2545_o;
  reg [9:0] n2546_o;
  reg n2547_o;
  wire [29:0] n2548_o;
  wire n2555_o;
  wire n2556_o;
  wire n2557_o;
  wire n2558_o;
  wire n2559_o;
  wire n2561_o;
  wire n2562_o;
  wire n2563_o;
  wire n2564_o;
  wire n2566_o;
  wire n2567_o;
  wire n2568_o;
  wire n2574_o;
  wire n2575_o;
  wire n2576_o;
  wire n2577_o;
  wire n2578_o;
  wire n2581_o;
  wire n2583_o;
  wire [20:0] n2586_o;
  reg [20:0] n2587_q;
  reg [1:0] n2588_q;
  reg [26:0] n2589_q;
  wire [29:0] n2590_o;
  reg n2591_q;
  reg [29:0] n2592_q;
  wire [30:0] n2593_o;
  wire [21:0] n2594_o;
  wire [21:0] n2595_o;
  reg [31:0] n2596_q;
  reg n2597_q;
  reg n2598_q;
  reg n2599_q;
  reg n2600_q;
  wire n2601_o;
  wire n2602_o;
  wire n2603_o;
  wire n2604_o;
  wire n2605_o;
  wire n2606_o;
  wire n2607_o;
  wire n2608_o;
  wire [1:0] n2609_o;
  reg n2610_o;
  wire [1:0] n2611_o;
  reg n2612_o;
  wire n2613_o;
  wire n2614_o;
  assign data_o = n2596_q;
  assign ack_o = n2597_q;
  assign clkgen_en_o = n2201_o;
  assign uart_txd_o = n2437_o;
  assign uart_rts_o = n2598_q;
  assign irq_rx_o = n2599_q;
  assign irq_tx_o = n2600_q;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:152:10  */
  assign acc_en = n2109_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:153:10  */
  assign addr = n2115_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:154:10  */
  assign wren = n2116_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:155:10  */
  assign rden = n2117_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:158:10  */
  assign uart_clk = n2614_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:173:10  */
  assign ctrl = n2587_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:185:10  */
  assign tx_engine = n2590_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:197:10  */
  assign rx_engine = n2593_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:210:10  */
  assign rx_fifo = n2594_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:210:19  */
  assign tx_fifo = n2595_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:226:29  */
  assign n2106_o = addr_i[8:3];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:226:56  */
  assign n2108_o = n2106_o == 6'b110100;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:226:17  */
  assign n2109_o = n2108_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:227:56  */
  assign n2111_o = addr_i[2];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:227:48  */
  assign n2113_o = {29'b11111111111111111111111110100, n2111_o};
  /* ../neorv32/rtl/core/neorv32_uart.vhd:227:78  */
  assign n2115_o = {n2113_o, 2'b00};
  /* ../neorv32/rtl/core/neorv32_uart.vhd:228:20  */
  assign n2116_o = acc_en & wren_i;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:229:20  */
  assign n2117_o = acc_en & rden_i;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:234:16  */
  assign n2119_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:247:18  */
  assign n2132_o = addr == 32'b11111111111111111111111110100000;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:248:39  */
  assign n2133_o = data_i[0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:249:39  */
  assign n2134_o = data_i[1];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:250:39  */
  assign n2135_o = data_i[2];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:251:39  */
  assign n2136_o = data_i[5:3];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:252:39  */
  assign n2137_o = data_i[15:6];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:254:39  */
  assign n2138_o = data_i[22];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:255:39  */
  assign n2139_o = data_i[23];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:256:39  */
  assign n2140_o = data_i[24];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:257:39  */
  assign n2141_o = data_i[25];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:258:39  */
  assign n2142_o = data_i[26];
  assign n2143_o = {n2142_o, n2141_o, n2140_o, n2139_o, n2138_o, n2137_o, n2136_o, n2135_o, n2134_o, n2133_o};
  /* ../neorv32/rtl/core/neorv32_uart.vhd:246:7  */
  assign n2145_o = wren & n2132_o;
  assign n2147_o = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 10'b0000000000, 3'b000, 1'b0, 1'b0, 1'b0};
  /* ../neorv32/rtl/core/neorv32_uart.vhd:268:22  */
  assign n2152_o = wren | rden;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:271:18  */
  assign n2154_o = addr == 32'b11111111111111111111111110100000;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:272:60  */
  assign n2155_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:273:60  */
  assign n2156_o = ctrl[1];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:274:60  */
  assign n2157_o = ctrl[2];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:275:60  */
  assign n2158_o = ctrl[5:3];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:276:60  */
  assign n2159_o = ctrl[15:6];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:278:63  */
  assign n2160_o = rx_fifo[20];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:279:63  */
  assign n2161_o = rx_fifo[21];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:280:67  */
  assign n2162_o = rx_fifo[19];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:280:55  */
  assign n2163_o = ~n2162_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:281:67  */
  assign n2164_o = tx_fifo[20];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:281:55  */
  assign n2165_o = ~n2164_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:282:67  */
  assign n2166_o = tx_fifo[21];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:282:55  */
  assign n2167_o = ~n2166_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:283:67  */
  assign n2168_o = tx_fifo[19];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:283:55  */
  assign n2169_o = ~n2168_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:285:60  */
  assign n2170_o = ctrl[16];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:286:60  */
  assign n2171_o = ctrl[17];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:287:60  */
  assign n2172_o = ctrl[18];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:288:60  */
  assign n2173_o = ctrl[19];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:289:60  */
  assign n2174_o = ctrl[20];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:291:65  */
  assign n2175_o = rx_engine[30];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:292:65  */
  assign n2176_o = tx_engine[27];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:292:81  */
  assign n2177_o = tx_fifo[20];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:292:70  */
  assign n2178_o = n2176_o | n2177_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:294:41  */
  assign n2179_o = rx_fifo[18:11];
  assign n2180_o = {n2174_o, n2173_o, n2172_o, n2171_o, n2170_o, n2169_o, n2167_o, n2165_o, n2163_o, n2161_o, n2160_o, n2159_o, n2158_o, n2157_o, n2156_o, n2155_o};
  assign n2181_o = {n2178_o, n2175_o};
  assign n2182_o = n2180_o[7:0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:271:9  */
  assign n2183_o = n2154_o ? n2182_o : n2179_o;
  assign n2184_o = n2180_o[26:8];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:271:9  */
  assign n2186_o = n2154_o ? n2184_o : 19'b0000000000000000000;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:271:9  */
  assign n2188_o = n2154_o ? n2181_o : 2'b00;
  assign n2189_o = {n2186_o, n2183_o};
  /* ../neorv32/rtl/core/neorv32_uart.vhd:270:7  */
  assign n2191_o = rden ? n2189_o : 27'b000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:270:7  */
  assign n2193_o = rden ? n2188_o : 2'b00;
  assign n2196_o = n2194_o[29:27];
  assign n2197_o = {n2193_o, n2196_o, n2191_o};
  /* ../neorv32/rtl/core/neorv32_uart.vhd:301:23  */
  assign n2201_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:302:52  */
  assign n2202_o = ctrl[5:3];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:320:24  */
  assign n2206_o = tx_fifo[0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:321:16  */
  assign tx_engine_fifo_inst_n2207 = tx_engine_fifo_inst_half_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:323:24  */
  assign n2208_o = tx_fifo[10:3];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:324:24  */
  assign n2209_o = tx_fifo[1];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:325:16  */
  assign tx_engine_fifo_inst_n2210 = tx_engine_fifo_inst_free_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:327:24  */
  assign n2211_o = tx_fifo[2];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:328:16  */
  assign tx_engine_fifo_inst_n2212 = tx_engine_fifo_inst_rdata_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:329:16  */
  assign tx_engine_fifo_inst_n2213 = tx_engine_fifo_inst_avail_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:309:3  */
  neorv32_fifo_256_8_9159cb8bcee7fcb95582f140960cdae72788d326 tx_engine_fifo_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .clear_i(n2206_o),
    .wdata_i(n2208_o),
    .we_i(n2209_o),
    .re_i(n2211_o),
    .half_o(tx_engine_fifo_inst_half_o),
    .free_o(tx_engine_fifo_inst_free_o),
    .rdata_o(tx_engine_fifo_inst_rdata_o),
    .avail_o(tx_engine_fifo_inst_avail_o));
  /* ../neorv32/rtl/core/neorv32_uart.vhd:332:35  */
  assign n2223_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:332:42  */
  assign n2224_o = ~n2223_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:332:58  */
  assign n2225_o = ctrl[1];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:332:49  */
  assign n2226_o = n2224_o | n2225_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:332:24  */
  assign n2227_o = n2226_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:333:26  */
  assign n2229_o = data_i[7:0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:334:52  */
  assign n2232_o = addr == 32'b11111111111111111111111110100100;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:334:42  */
  assign n2233_o = wren & n2232_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:334:24  */
  assign n2234_o = n2233_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:335:40  */
  assign n2237_o = tx_engine[2:0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:335:46  */
  assign n2239_o = n2237_o == 3'b100;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:335:24  */
  assign n2240_o = n2239_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:341:24  */
  assign n2244_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:342:25  */
  assign n2245_o = ctrl[19];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:342:55  */
  assign n2246_o = tx_fifo[20];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:342:43  */
  assign n2247_o = ~n2246_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:342:38  */
  assign n2248_o = n2245_o & n2247_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:343:25  */
  assign n2249_o = ctrl[20];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:343:55  */
  assign n2250_o = tx_fifo[21];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:343:43  */
  assign n2251_o = ~n2250_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:343:38  */
  assign n2252_o = n2249_o & n2251_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:342:63  */
  assign n2253_o = n2248_o | n2252_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:341:31  */
  assign n2254_o = n2244_o & n2253_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:360:24  */
  assign n2257_o = rx_fifo[0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:361:16  */
  assign rx_engine_fifo_inst_n2258 = rx_engine_fifo_inst_half_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:363:24  */
  assign n2259_o = rx_fifo[10:3];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:364:24  */
  assign n2260_o = rx_fifo[1];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:365:16  */
  assign rx_engine_fifo_inst_n2261 = rx_engine_fifo_inst_free_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:367:24  */
  assign n2262_o = rx_fifo[2];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:368:16  */
  assign rx_engine_fifo_inst_n2263 = rx_engine_fifo_inst_rdata_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:369:16  */
  assign rx_engine_fifo_inst_n2264 = rx_engine_fifo_inst_avail_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_uart.vhd:349:3  */
  neorv32_fifo_256_8_9159cb8bcee7fcb95582f140960cdae72788d326 rx_engine_fifo_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .clear_i(n2257_o),
    .wdata_i(n2259_o),
    .we_i(n2260_o),
    .re_i(n2262_o),
    .half_o(rx_engine_fifo_inst_half_o),
    .free_o(rx_engine_fifo_inst_free_o),
    .rdata_o(rx_engine_fifo_inst_rdata_o),
    .avail_o(rx_engine_fifo_inst_avail_o));
  /* ../neorv32/rtl/core/neorv32_uart.vhd:372:35  */
  assign n2274_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:372:42  */
  assign n2275_o = ~n2274_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:372:58  */
  assign n2276_o = ctrl[1];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:372:49  */
  assign n2277_o = n2275_o | n2276_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:372:24  */
  assign n2278_o = n2277_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:373:34  */
  assign n2280_o = rx_engine[10:3];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:374:30  */
  assign n2281_o = rx_engine[26];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:375:52  */
  assign n2284_o = addr == 32'b11111111111111111111111110100100;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:375:42  */
  assign n2285_o = rden & n2284_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:375:24  */
  assign n2286_o = n2285_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:381:24  */
  assign n2290_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:382:25  */
  assign n2291_o = ctrl[16];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:382:51  */
  assign n2292_o = rx_fifo[20];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:382:39  */
  assign n2293_o = n2291_o & n2292_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:383:25  */
  assign n2294_o = ctrl[17];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:383:51  */
  assign n2295_o = rx_fifo[21];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:383:39  */
  assign n2296_o = n2294_o & n2295_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:382:58  */
  assign n2297_o = n2293_o | n2296_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:384:25  */
  assign n2298_o = ctrl[18];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:384:56  */
  assign n2299_o = rx_fifo[19];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:384:44  */
  assign n2300_o = ~n2299_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:384:39  */
  assign n2301_o = n2298_o & n2300_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:383:58  */
  assign n2302_o = n2297_o | n2301_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:381:31  */
  assign n2303_o = n2290_o & n2302_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:395:47  */
  assign n2308_o = tx_engine[28];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:395:51  */
  assign n2309_o = {n2308_o, uart_cts_i};
  /* ../neorv32/rtl/core/neorv32_uart.vhd:401:34  */
  assign n2311_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:402:22  */
  assign n2312_o = tx_engine[2:0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:406:37  */
  assign n2313_o = ctrl[15:6];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:408:40  */
  assign n2315_o = tx_fifo[18:11];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:408:46  */
  assign n2317_o = {n2315_o, 1'b0};
  /* ../neorv32/rtl/core/neorv32_uart.vhd:409:23  */
  assign n2318_o = tx_fifo[20];
  assign n2320_o = tx_engine[1:0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:409:11  */
  assign n2321_o = n2318_o ? 2'b01 : n2320_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:404:9  */
  assign n2323_o = n2312_o == 3'b100;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:415:33  */
  assign n2324_o = tx_engine[29];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:415:37  */
  assign n2325_o = ~n2324_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:415:53  */
  assign n2326_o = ctrl[2];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:415:61  */
  assign n2327_o = ~n2326_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:415:44  */
  assign n2328_o = n2325_o | n2327_o;
  assign n2330_o = tx_engine[1:0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:415:11  */
  assign n2331_o = n2328_o ? 2'b11 : n2330_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:413:9  */
  assign n2333_o = n2312_o == 3'b101;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:422:39  */
  assign n2335_o = tx_engine[25:16];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2341_o = n2335_o[9];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2343_o = 1'b0 | n2341_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2345_o = n2335_o[8];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2346_o = n2343_o | n2345_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2347_o = n2335_o[7];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2348_o = n2346_o | n2347_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2349_o = n2335_o[6];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2350_o = n2348_o | n2349_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2351_o = n2335_o[5];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2352_o = n2350_o | n2351_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2353_o = n2335_o[4];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2354_o = n2352_o | n2353_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2355_o = n2335_o[3];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2356_o = n2354_o | n2355_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2357_o = n2335_o[2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2358_o = n2356_o | n2357_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2359_o = n2335_o[1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2360_o = n2358_o | n2359_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2361_o = n2335_o[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2362_o = n2360_o | n2361_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:422:48  */
  assign n2363_o = ~n2362_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:423:41  */
  assign n2364_o = ctrl[15:6];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:424:73  */
  assign n2365_o = tx_engine[15:12];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:424:81  */
  assign n2367_o = n2365_o - 4'b0001;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:425:56  */
  assign n2368_o = tx_engine[11:4];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:425:40  */
  assign n2370_o = {1'b1, n2368_o};
  /* ../neorv32/rtl/core/neorv32_uart.vhd:427:73  */
  assign n2371_o = tx_engine[25:16];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:427:82  */
  assign n2373_o = n2371_o - 10'b0000000001;
  assign n2374_o = {n2364_o, n2367_o, n2370_o};
  assign n2375_o = n2374_o[12:0];
  assign n2376_o = tx_engine[15:3];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:422:13  */
  assign n2377_o = n2363_o ? n2375_o : n2376_o;
  assign n2378_o = n2374_o[22:13];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:422:13  */
  assign n2379_o = n2363_o ? n2378_o : n2373_o;
  assign n2380_o = {n2379_o, n2377_o};
  assign n2381_o = tx_engine[25:3];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:421:11  */
  assign n2382_o = uart_clk ? n2380_o : n2381_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:430:37  */
  assign n2384_o = tx_engine[15:12];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2390_o = n2384_o[3];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2392_o = 1'b0 | n2390_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2394_o = n2384_o[2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2395_o = n2392_o | n2394_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2396_o = n2384_o[1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2397_o = n2395_o | n2396_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2398_o = n2384_o[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2399_o = n2397_o | n2398_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:430:45  */
  assign n2400_o = ~n2399_o;
  assign n2403_o = tx_engine[1:0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:430:11  */
  assign n2404_o = n2400_o ? 2'b00 : n2403_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:430:11  */
  assign n2405_o = n2400_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:419:9  */
  assign n2407_o = n2312_o == 3'b111;
  assign n2409_o = {n2407_o, n2333_o, n2323_o};
  /* ../neorv32/rtl/core/neorv32_uart.vhd:402:7  */
  always @*
    case (n2409_o)
      3'b100: n2410_o = n2404_o;
      3'b010: n2410_o = n2331_o;
      3'b001: n2410_o = n2321_o;
      default: n2410_o = 2'b00;
    endcase
  assign n2411_o = n2382_o[8:0];
  assign n2412_o = tx_engine[11:3];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:402:7  */
  always @*
    case (n2409_o)
      3'b100: n2413_o = n2411_o;
      3'b010: n2413_o = n2412_o;
      3'b001: n2413_o = n2317_o;
      default: n2413_o = n2412_o;
    endcase
  assign n2414_o = n2382_o[12:9];
  assign n2415_o = tx_engine[15:12];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:402:7  */
  always @*
    case (n2409_o)
      3'b100: n2416_o = n2414_o;
      3'b010: n2416_o = n2415_o;
      3'b001: n2416_o = 4'b1011;
      default: n2416_o = n2415_o;
    endcase
  assign n2417_o = n2382_o[22:13];
  assign n2418_o = tx_engine[25:16];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:402:7  */
  always @*
    case (n2409_o)
      3'b100: n2419_o = n2417_o;
      3'b010: n2419_o = n2418_o;
      3'b001: n2419_o = n2313_o;
      default: n2419_o = n2418_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_uart.vhd:402:7  */
  always @*
    case (n2409_o)
      3'b100: n2420_o = n2405_o;
      3'b010: n2420_o = 1'b0;
      3'b001: n2420_o = 1'b0;
      default: n2420_o = 1'b0;
    endcase
  assign n2421_o = {n2420_o, n2419_o, n2416_o, n2413_o, n2311_o, n2410_o};
  /* ../neorv32/rtl/core/neorv32_uart.vhd:444:46  */
  assign n2428_o = tx_engine[1:0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:444:59  */
  assign n2430_o = n2428_o == 2'b00;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:444:25  */
  assign n2431_o = n2430_o ? 1'b0 : 1'b1;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:447:31  */
  assign n2433_o = tx_engine[3];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:447:51  */
  assign n2434_o = tx_engine[2:0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:447:57  */
  assign n2436_o = n2434_o == 3'b111;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:447:35  */
  assign n2437_o = n2436_o ? n2433_o : 1'b1;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:458:44  */
  assign n2441_o = rx_engine[29];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:459:44  */
  assign n2442_o = rx_engine[28];
  assign n2443_o = {n2441_o, n2442_o};
  assign n2444_o = rx_engine[28:27];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:457:7  */
  assign n2445_o = uart_clk ? n2443_o : n2444_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:466:34  */
  assign n2447_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:467:22  */
  assign n2448_o = rx_engine[1:0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:471:47  */
  assign n2449_o = ctrl[15:7];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:471:36  */
  assign n2451_o = {1'b0, n2449_o};
  /* ../neorv32/rtl/core/neorv32_uart.vhd:473:29  */
  assign n2453_o = rx_engine[28:27];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:473:42  */
  assign n2455_o = n2453_o == 2'b01;
  assign n2457_o = rx_engine[0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:473:11  */
  assign n2458_o = n2455_o ? 1'b1 : n2457_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:469:9  */
  assign n2460_o = n2448_o == 2'b10;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:480:39  */
  assign n2462_o = rx_engine[25:16];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2468_o = n2462_o[9];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2470_o = 1'b0 | n2468_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2472_o = n2462_o[8];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2473_o = n2470_o | n2472_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2474_o = n2462_o[7];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2475_o = n2473_o | n2474_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2476_o = n2462_o[6];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2477_o = n2475_o | n2476_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2478_o = n2462_o[5];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2479_o = n2477_o | n2478_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2480_o = n2462_o[4];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2481_o = n2479_o | n2480_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2482_o = n2462_o[3];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2483_o = n2481_o | n2482_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2484_o = n2462_o[2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2485_o = n2483_o | n2484_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2486_o = n2462_o[1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2487_o = n2485_o | n2486_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2488_o = n2462_o[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2489_o = n2487_o | n2488_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:480:48  */
  assign n2490_o = ~n2489_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:481:41  */
  assign n2491_o = ctrl[15:6];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:482:73  */
  assign n2492_o = rx_engine[15:12];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:482:81  */
  assign n2494_o = n2492_o - 4'b0001;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:483:50  */
  assign n2495_o = rx_engine[29];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:483:70  */
  assign n2496_o = rx_engine[11:3];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:483:54  */
  assign n2497_o = {n2495_o, n2496_o};
  /* ../neorv32/rtl/core/neorv32_uart.vhd:485:73  */
  assign n2498_o = rx_engine[25:16];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:485:82  */
  assign n2500_o = n2498_o - 10'b0000000001;
  assign n2501_o = {n2491_o, n2494_o, n2497_o};
  assign n2502_o = n2501_o[13:0];
  assign n2503_o = rx_engine[15:2];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:480:13  */
  assign n2504_o = n2490_o ? n2502_o : n2503_o;
  assign n2505_o = n2501_o[23:14];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:480:13  */
  assign n2506_o = n2490_o ? n2505_o : n2500_o;
  assign n2507_o = {n2506_o, n2504_o};
  assign n2508_o = rx_engine[25:2];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:479:11  */
  assign n2509_o = uart_clk ? n2507_o : n2508_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:488:37  */
  assign n2511_o = rx_engine[15:12];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2517_o = n2511_o[3];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2519_o = 1'b0 | n2517_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2521_o = n2511_o[2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2522_o = n2519_o | n2521_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2523_o = n2511_o[1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2524_o = n2522_o | n2523_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n2525_o = n2511_o[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n2526_o = n2524_o | n2525_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:488:45  */
  assign n2527_o = ~n2526_o;
  assign n2530_o = rx_engine[0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:488:11  */
  assign n2531_o = n2527_o ? 1'b0 : n2530_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:488:11  */
  assign n2532_o = n2527_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:477:9  */
  assign n2534_o = n2448_o == 2'b11;
  assign n2536_o = {n2534_o, n2460_o};
  /* ../neorv32/rtl/core/neorv32_uart.vhd:467:7  */
  always @*
    case (n2536_o)
      2'b10: n2537_o = n2531_o;
      2'b01: n2537_o = n2458_o;
      default: n2537_o = 1'b0;
    endcase
  assign n2538_o = n2509_o[9:0];
  assign n2539_o = rx_engine[11:2];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:467:7  */
  always @*
    case (n2536_o)
      2'b10: n2540_o = n2538_o;
      2'b01: n2540_o = n2539_o;
      default: n2540_o = n2539_o;
    endcase
  assign n2541_o = n2509_o[13:10];
  assign n2542_o = rx_engine[15:12];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:467:7  */
  always @*
    case (n2536_o)
      2'b10: n2543_o = n2541_o;
      2'b01: n2543_o = 4'b1010;
      default: n2543_o = n2542_o;
    endcase
  assign n2544_o = n2509_o[23:14];
  assign n2545_o = rx_engine[25:16];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:467:7  */
  always @*
    case (n2536_o)
      2'b10: n2546_o = n2544_o;
      2'b01: n2546_o = n2451_o;
      default: n2546_o = n2545_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_uart.vhd:467:7  */
  always @*
    case (n2536_o)
      2'b10: n2547_o = n2532_o;
      2'b01: n2547_o = 1'b0;
      default: n2547_o = 1'b0;
    endcase
  assign n2548_o = {uart_rxd_i, n2445_o, n2547_o, n2546_o, n2543_o, n2540_o, n2447_o, n2537_o};
  /* ../neorv32/rtl/core/neorv32_uart.vhd:505:34  */
  assign n2555_o = addr == 32'b11111111111111111111111110100100;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:505:24  */
  assign n2556_o = rden & n2555_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:505:66  */
  assign n2557_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:505:73  */
  assign n2558_o = ~n2557_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:505:57  */
  assign n2559_o = n2556_o | n2558_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:507:22  */
  assign n2561_o = rx_fifo[1];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:507:45  */
  assign n2562_o = rx_fifo[19];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:507:50  */
  assign n2563_o = ~n2562_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:507:32  */
  assign n2564_o = n2561_o & n2563_o;
  assign n2566_o = rx_engine[30];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:507:7  */
  assign n2567_o = n2564_o ? 1'b1 : n2566_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:505:7  */
  assign n2568_o = n2559_o ? 1'b0 : n2567_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:517:16  */
  assign n2574_o = ctrl[2];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:518:18  */
  assign n2575_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:518:25  */
  assign n2576_o = ~n2575_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:519:21  */
  assign n2577_o = rx_fifo[21];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:518:32  */
  assign n2578_o = n2576_o | n2577_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:518:9  */
  assign n2581_o = n2578_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:517:7  */
  assign n2583_o = n2574_o ? n2581_o : 1'b0;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:245:5  */
  assign n2586_o = n2145_o ? n2143_o : ctrl;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:245:5  */
  always @(posedge clk_i or posedge n2119_o)
    if (n2119_o)
      n2587_q <= n2147_o;
    else
      n2587_q <= n2586_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:393:5  */
  always @(posedge clk_i)
    n2588_q <= n2309_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:393:5  */
  always @(posedge clk_i)
    n2589_q <= n2421_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:393:5  */
  assign n2590_o = {n2588_q, n2431_o, n2589_q};
  /* ../neorv32/rtl/core/neorv32_uart.vhd:504:5  */
  always @(posedge clk_i)
    n2591_q <= n2568_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:454:5  */
  always @(posedge clk_i)
    n2592_q <= n2548_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:454:5  */
  assign n2593_o = {n2591_q, n2592_q};
  assign n2594_o = {rx_engine_fifo_inst_n2258, rx_engine_fifo_inst_n2264, rx_engine_fifo_inst_n2261, rx_engine_fifo_inst_n2263, n2280_o, n2286_o, n2281_o, n2278_o};
  assign n2595_o = {tx_engine_fifo_inst_n2207, tx_engine_fifo_inst_n2213, tx_engine_fifo_inst_n2210, tx_engine_fifo_inst_n2212, n2229_o, n2240_o, n2234_o, n2227_o};
  /* ../neorv32/rtl/core/neorv32_uart.vhd:267:5  */
  always @(posedge clk_i)
    n2596_q <= n2197_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:267:5  */
  always @(posedge clk_i)
    n2597_q <= n2152_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:516:5  */
  always @(posedge clk_i)
    n2598_q <= n2583_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:380:5  */
  always @(posedge clk_i)
    n2599_q <= n2303_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:340:5  */
  always @(posedge clk_i)
    n2600_q <= n2254_o;
  /* ../neorv32/rtl/core/neorv32_uart.vhd:369:16  */
  assign n2601_o = clkgen_i[0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:368:16  */
  assign n2602_o = clkgen_i[1];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:365:16  */
  assign n2603_o = clkgen_i[2];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:361:16  */
  assign n2604_o = clkgen_i[3];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:349:3  */
  assign n2605_o = clkgen_i[4];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:349:3  */
  assign n2606_o = clkgen_i[5];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:349:3  */
  assign n2607_o = clkgen_i[6];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:349:3  */
  assign n2608_o = clkgen_i[7];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:302:26  */
  assign n2609_o = n2202_o[1:0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:302:26  */
  always @*
    case (n2609_o)
      2'b00: n2610_o = n2601_o;
      2'b01: n2610_o = n2602_o;
      2'b10: n2610_o = n2603_o;
      2'b11: n2610_o = n2604_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_uart.vhd:302:26  */
  assign n2611_o = n2202_o[1:0];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:302:26  */
  always @*
    case (n2611_o)
      2'b00: n2612_o = n2605_o;
      2'b01: n2612_o = n2606_o;
      2'b10: n2612_o = n2607_o;
      2'b11: n2612_o = n2608_o;
    endcase
  /* ../neorv32/rtl/core/neorv32_uart.vhd:302:26  */
  assign n2613_o = n2202_o[2];
  /* ../neorv32/rtl/core/neorv32_uart.vhd:302:26  */
  assign n2614_o = n2613_o ? n2612_o : n2610_o;
endmodule

module neorv32_mtime
  (input  clk_i,
   input  rstn_i,
   input  [31:0] addr_i,
   input  rden_i,
   input  wren_i,
   input  [31:0] data_i,
   output [31:0] data_o,
   output ack_o,
   output irq_o);
  wire acc_en;
  wire [31:0] addr;
  wire wren;
  wire rden;
  wire mtime_lo_we;
  wire mtime_hi_we;
  wire [31:0] mtimecmp_lo;
  wire [31:0] mtimecmp_hi;
  wire [31:0] mtime_lo;
  wire [32:0] mtime_lo_nxt;
  wire mtime_lo_ovfl;
  wire [31:0] mtime_hi;
  wire cmp_lo_ge;
  wire cmp_lo_ge_ff;
  wire cmp_hi_eq;
  wire cmp_hi_gt;
  wire [4:0] n1977_o;
  wire n1979_o;
  wire n1980_o;
  wire [1:0] n1982_o;
  wire [29:0] n1984_o;
  wire [31:0] n1986_o;
  wire n1987_o;
  wire n1988_o;
  wire n1990_o;
  wire n1993_o;
  wire n1996_o;
  wire n1998_o;
  wire n1999_o;
  wire n2001_o;
  wire n2002_o;
  wire n2005_o;
  wire n2008_o;
  wire n2009_o;
  wire n2012_o;
  wire [31:0] n2014_o;
  wire [31:0] n2015_o;
  wire n2016_o;
  wire [31:0] n2017_o;
  wire [31:0] n2018_o;
  wire [31:0] n2019_o;
  wire [32:0] n2043_o;
  wire [32:0] n2045_o;
  wire n2048_o;
  wire [1:0] n2049_o;
  wire n2051_o;
  wire n2053_o;
  wire n2055_o;
  wire [2:0] n2056_o;
  reg [31:0] n2057_o;
  wire [31:0] n2059_o;
  wire n2066_o;
  wire n2067_o;
  wire n2072_o;
  wire n2073_o;
  wire n2076_o;
  wire n2077_o;
  wire n2080_o;
  wire n2081_o;
  reg n2083_q;
  reg n2084_q;
  wire [31:0] n2085_o;
  reg [31:0] n2086_q;
  wire [31:0] n2087_o;
  reg [31:0] n2088_q;
  reg [31:0] n2089_q;
  reg n2090_q;
  reg [31:0] n2091_q;
  reg n2092_q;
  reg [31:0] n2093_q;
  reg n2094_q;
  reg n2095_q;
  assign data_o = n2093_q;
  assign ack_o = n2094_q;
  assign irq_o = n2095_q;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:68:10  */
  assign acc_en = n1980_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:69:10  */
  assign addr = n1986_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:70:10  */
  assign wren = n1987_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:71:10  */
  assign rden = n1988_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:74:10  */
  assign mtime_lo_we = n2083_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:75:10  */
  assign mtime_hi_we = n2084_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:78:10  */
  assign mtimecmp_lo = n2086_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:79:10  */
  assign mtimecmp_hi = n2088_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:80:10  */
  assign mtime_lo = n2089_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:81:10  */
  assign mtime_lo_nxt = n2045_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:82:10  */
  assign mtime_lo_ovfl = n2090_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:83:10  */
  assign mtime_hi = n2091_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:86:10  */
  assign cmp_lo_ge = n2073_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:87:10  */
  assign cmp_lo_ge_ff = n2092_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:88:10  */
  assign cmp_hi_eq = n2077_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:89:10  */
  assign cmp_hi_gt = n2081_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:95:29  */
  assign n1977_o = addr_i[8:4];
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:95:56  */
  assign n1979_o = n1977_o == 5'b11001;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:95:17  */
  assign n1980_o = n1979_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:96:54  */
  assign n1982_o = addr_i[3:2];
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:96:46  */
  assign n1984_o = {28'b1111111111111111111111111001, n1982_o};
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:96:76  */
  assign n1986_o = {n1984_o, 2'b00};
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:97:20  */
  assign n1987_o = acc_en & wren_i;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:98:20  */
  assign n1988_o = acc_en & rden_i;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:105:16  */
  assign n1990_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:116:18  */
  assign n1993_o = addr == 32'b11111111111111111111111110011000;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:119:18  */
  assign n1996_o = addr == 32'b11111111111111111111111110011100;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:115:7  */
  assign n1998_o = wren & n1993_o;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:115:7  */
  assign n1999_o = wren & n1996_o;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:126:33  */
  assign n2001_o = addr == 32'b11111111111111111111111110010000;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:126:23  */
  assign n2002_o = wren & n2001_o;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:126:7  */
  assign n2005_o = n2002_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:131:33  */
  assign n2008_o = addr == 32'b11111111111111111111111110010100;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:131:23  */
  assign n2009_o = wren & n2008_o;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:131:7  */
  assign n2012_o = n2009_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:139:33  */
  assign n2014_o = mtime_lo_nxt[31:0];
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:136:7  */
  assign n2015_o = mtime_lo_we ? data_i : n2014_o;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:141:39  */
  assign n2016_o = mtime_lo_nxt[32];
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:147:58  */
  assign n2017_o = {31'b0, mtime_lo_ovfl};  //  uext
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:147:58  */
  assign n2018_o = mtime_hi + n2017_o;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:144:7  */
  assign n2019_o = mtime_hi_we ? data_i : n2018_o;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:153:50  */
  assign n2043_o = {1'b0, mtime_lo};
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:153:62  */
  assign n2045_o = n2043_o + 33'b000000000000000000000000000000001;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:161:22  */
  assign n2048_o = rden | wren;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:164:18  */
  assign n2049_o = addr[3:2];
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:165:11  */
  assign n2051_o = n2049_o == 2'b00;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:166:11  */
  assign n2053_o = n2049_o == 2'b01;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:167:11  */
  assign n2055_o = n2049_o == 2'b10;
  assign n2056_o = {n2055_o, n2053_o, n2051_o};
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:164:9  */
  always @*
    case (n2056_o)
      3'b100: n2057_o = mtimecmp_lo;
      3'b010: n2057_o = mtime_hi;
      3'b001: n2057_o = mtime_lo;
      default: n2057_o = mtimecmp_hi;
    endcase
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:163:7  */
  assign n2059_o = rden ? n2057_o : 32'b00000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:181:47  */
  assign n2066_o = cmp_hi_eq & cmp_lo_ge_ff;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:181:33  */
  assign n2067_o = cmp_hi_gt | n2066_o;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:186:45  */
  assign n2072_o = $unsigned(mtime_lo) >= $unsigned(mtimecmp_lo);
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:186:20  */
  assign n2073_o = n2072_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:187:45  */
  assign n2076_o = mtime_hi == mtimecmp_hi;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:187:20  */
  assign n2077_o = n2076_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:188:45  */
  assign n2080_o = $unsigned(mtime_hi) > $unsigned(mtimecmp_hi);
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:188:20  */
  assign n2081_o = n2080_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:113:5  */
  always @(posedge clk_i or posedge n1990_o)
    if (n1990_o)
      n2083_q <= 1'b0;
    else
      n2083_q <= n2005_o;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:113:5  */
  always @(posedge clk_i or posedge n1990_o)
    if (n1990_o)
      n2084_q <= 1'b0;
    else
      n2084_q <= n2012_o;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:113:5  */
  assign n2085_o = n1998_o ? data_i : mtimecmp_lo;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:113:5  */
  always @(posedge clk_i or posedge n1990_o)
    if (n1990_o)
      n2086_q <= 32'b00000000000000000000000000000000;
    else
      n2086_q <= n2085_o;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:113:5  */
  assign n2087_o = n1999_o ? data_i : mtimecmp_hi;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:113:5  */
  always @(posedge clk_i or posedge n1990_o)
    if (n1990_o)
      n2088_q <= 32'b00000000000000000000000000000000;
    else
      n2088_q <= n2087_o;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:113:5  */
  always @(posedge clk_i or posedge n1990_o)
    if (n1990_o)
      n2089_q <= 32'b00000000000000000000000000000000;
    else
      n2089_q <= n2015_o;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:113:5  */
  always @(posedge clk_i or posedge n1990_o)
    if (n1990_o)
      n2090_q <= 1'b0;
    else
      n2090_q <= n2016_o;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:113:5  */
  always @(posedge clk_i or posedge n1990_o)
    if (n1990_o)
      n2091_q <= 32'b00000000000000000000000000000000;
    else
      n2091_q <= n2019_o;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:179:5  */
  always @(posedge clk_i)
    n2092_q <= cmp_lo_ge;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:160:5  */
  always @(posedge clk_i)
    n2093_q <= n2059_o;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:160:5  */
  always @(posedge clk_i)
    n2094_q <= n2048_o;
  /* ../neorv32/rtl/core/neorv32_mtime.vhd:179:5  */
  always @(posedge clk_i)
    n2095_q <= n2067_o;
endmodule

module neorv32_wishbone_1024_2048_255_faf1cd4bdf2d59261beed066baf3c3e69ee5d9f7
  (input  clk_i,
   input  rstn_i,
   input  src_i,
   input  [31:0] addr_i,
   input  rden_i,
   input  wren_i,
   input  [3:0] ben_i,
   input  [31:0] data_i,
   input  priv_i,
   input  xip_en_i,
   input  [3:0] xip_page_i,
   input  [31:0] wb_dat_i,
   input  wb_ack_i,
   input  wb_err_i,
   output [31:0] data_o,
   output ack_o,
   output err_o,
   output tmo_o,
   output ext_o,
   output [2:0] wb_tag_o,
   output [31:0] wb_adr_o,
   output [31:0] wb_dat_o,
   output wb_we_o,
   output [3:0] wb_sel_o,
   output wb_stb_o,
   output wb_cyc_o);
  wire int_imem_acc;
  wire int_dmem_acc;
  wire int_boot_acc;
  wire xip_acc;
  wire xbus_access;
  wire [116:0] ctrl;
  wire stb_int;
  wire cyc_int;
  wire [31:0] rdata;
  wire [31:0] end_wdata;
  wire [3:0] end_byteen;
  wire ack_gated;
  wire [31:0] rdata_gated;
  wire [21:0] n1725_o;
  wire n1728_o;
  wire n1730_o;
  wire n1731_o;
  wire [20:0] n1735_o;
  wire n1738_o;
  wire n1740_o;
  wire n1741_o;
  wire [15:0] n1744_o;
  wire n1746_o;
  wire n1747_o;
  wire [3:0] n1750_o;
  wire n1751_o;
  wire n1752_o;
  wire n1753_o;
  wire n1755_o;
  wire n1756_o;
  wire n1757_o;
  wire n1758_o;
  wire n1759_o;
  wire n1760_o;
  wire n1761_o;
  wire n1763_o;
  wire n1778_o;
  wire n1785_o;
  wire n1786_o;
  wire n1787_o;
  wire n1788_o;
  wire [64:0] n1790_o;
  wire [1:0] n1791_o;
  wire n1792_o;
  wire n1793_o;
  wire [64:0] n1794_o;
  wire [64:0] n1795_o;
  wire [3:0] n1796_o;
  wire [3:0] n1797_o;
  wire [1:0] n1798_o;
  wire [1:0] n1799_o;
  wire [8:0] n1803_o;
  wire n1809_o;
  wire n1811_o;
  wire n1813_o;
  wire n1814_o;
  wire n1815_o;
  wire n1816_o;
  wire n1817_o;
  wire n1818_o;
  wire n1819_o;
  wire n1820_o;
  wire n1821_o;
  wire n1822_o;
  wire n1823_o;
  wire n1824_o;
  wire n1825_o;
  wire n1826_o;
  wire n1827_o;
  wire n1828_o;
  wire n1829_o;
  wire n1831_o;
  wire n1836_o;
  wire n1837_o;
  wire n1838_o;
  wire n1839_o;
  wire n1840_o;
  wire n1841_o;
  wire n1842_o;
  wire n1843_o;
  wire n1844_o;
  wire n1845_o;
  wire [8:0] n1846_o;
  wire [8:0] n1848_o;
  wire [11:0] n1849_o;
  wire n1850_o;
  wire n1852_o;
  wire [31:0] n1853_o;
  wire n1855_o;
  wire [11:0] n1856_o;
  wire [11:0] n1857_o;
  wire n1859_o;
  wire [116:0] n1860_o;
  wire [116:0] n1862_o;
  wire n1865_o;
  wire [7:0] n1872_o;
  wire [7:0] n1875_o;
  wire [7:0] n1877_o;
  wire [7:0] n1879_o;
  wire [31:0] n1880_o;
  wire [31:0] n1882_o;
  wire n1889_o;
  wire n1892_o;
  wire n1894_o;
  wire n1896_o;
  wire [3:0] n1897_o;
  wire [3:0] n1899_o;
  wire n1900_o;
  wire n1901_o;
  wire n1903_o;
  wire [31:0] n1904_o;
  wire [31:0] n1906_o;
  wire [31:0] n1908_o;
  wire [31:0] n1910_o;
  wire [7:0] n1917_o;
  wire [7:0] n1920_o;
  wire [7:0] n1922_o;
  wire [7:0] n1924_o;
  wire [31:0] n1925_o;
  wire n1926_o;
  wire n1928_o;
  wire n1929_o;
  wire n1930_o;
  wire n1932_o;
  wire n1933_o;
  wire n1936_o;
  wire n1937_o;
  wire n1938_o;
  wire n1939_o;
  wire n1941_o;
  wire n1942_o;
  wire n1943_o;
  wire n1944_o;
  wire n1945_o;
  wire n1946_o;
  wire n1947_o;
  wire n1948_o;
  wire n1949_o;
  wire n1951_o;
  wire n1952_o;
  wire [31:0] n1954_o;
  wire [31:0] n1955_o;
  wire [31:0] n1957_o;
  wire [31:0] n1958_o;
  wire n1959_o;
  wire n1960_o;
  wire n1961_o;
  wire n1962_o;
  wire n1964_o;
  wire n1965_o;
  wire [3:0] n1967_o;
  wire [3:0] n1968_o;
  wire n1970_o;
  reg [116:0] n1971_q;
  wire [2:0] n1972_o;
  assign data_o = n1910_o;
  assign ack_o = n1928_o;
  assign err_o = n1929_o;
  assign tmo_o = n1930_o;
  assign ext_o = n1865_o;
  assign wb_tag_o = n1972_o;
  assign wb_adr_o = n1954_o;
  assign wb_dat_o = n1957_o;
  assign wb_we_o = n1964_o;
  assign wb_sel_o = n1967_o;
  assign wb_stb_o = n1970_o;
  assign wb_cyc_o = cyc_int;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:110:10  */
  assign int_imem_acc = n1731_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:111:10  */
  assign int_dmem_acc = n1741_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:112:10  */
  assign int_boot_acc = n1747_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:113:10  */
  assign xip_acc = n1753_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:114:10  */
  assign xbus_access = n1761_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:132:10  */
  assign ctrl = n1971_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:133:10  */
  assign stb_int = n1941_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:134:10  */
  assign cyc_int = n1951_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:135:10  */
  assign rdata = n1908_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:138:10  */
  assign end_wdata = n1882_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:139:10  */
  assign end_byteen = n1899_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:142:10  */
  assign ack_gated = n1901_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:143:10  */
  assign rdata_gated = n1904_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:166:35  */
  assign n1725_o = addr_i[31:10];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:166:79  */
  assign n1728_o = n1725_o == 22'b0000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:166:137  */
  assign n1730_o = n1728_o & 1'b1;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:166:23  */
  assign n1731_o = n1730_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:167:35  */
  assign n1735_o = addr_i[31:11];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:167:79  */
  assign n1738_o = n1735_o == 21'b100000000000000000000;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:167:137  */
  assign n1740_o = n1738_o & 1'b1;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:167:23  */
  assign n1741_o = n1740_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:169:35  */
  assign n1744_o = addr_i[31:16];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:169:50  */
  assign n1746_o = n1744_o == 16'b1111111111111111;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:169:23  */
  assign n1747_o = n1746_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:171:56  */
  assign n1750_o = addr_i[31:28];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:171:71  */
  assign n1751_o = n1750_o == xip_page_i;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:171:45  */
  assign n1752_o = xip_en_i & n1751_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:171:23  */
  assign n1753_o = n1752_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:173:20  */
  assign n1755_o = ~int_imem_acc;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:173:43  */
  assign n1756_o = ~int_dmem_acc;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:173:38  */
  assign n1757_o = n1755_o & n1756_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:173:66  */
  assign n1758_o = ~int_boot_acc;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:173:61  */
  assign n1759_o = n1757_o & n1758_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:173:89  */
  assign n1760_o = ~xip_acc;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:173:84  */
  assign n1761_o = n1759_o & n1760_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:180:16  */
  assign n1763_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:196:29  */
  assign n1778_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:204:16  */
  assign n1785_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:204:22  */
  assign n1786_o = ~n1785_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:206:45  */
  assign n1787_o = wren_i | rden_i;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:206:32  */
  assign n1788_o = xbus_access & n1787_o;
  assign n1790_o = {end_wdata, addr_i, wren_i};
  assign n1791_o = {priv_i, src_i};
  assign n1792_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:206:9  */
  assign n1793_o = n1788_o ? 1'b1 : n1792_o;
  assign n1794_o = ctrl[66:2];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:204:7  */
  assign n1795_o = n1852_o ? n1790_o : n1794_o;
  assign n1796_o = ctrl[102:99];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:204:7  */
  assign n1797_o = n1855_o ? end_byteen : n1796_o;
  assign n1798_o = ctrl[116:115];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:204:7  */
  assign n1799_o = n1859_o ? n1791_o : n1798_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:223:59  */
  assign n1803_o = ctrl[114:106];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n1809_o = n1803_o[8];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n1811_o = 1'b0 | n1809_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n1813_o = n1803_o[7];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n1814_o = n1811_o | n1813_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n1815_o = n1803_o[6];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n1816_o = n1814_o | n1815_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n1817_o = n1803_o[5];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n1818_o = n1816_o | n1817_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n1819_o = n1803_o[4];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n1820_o = n1818_o | n1819_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n1821_o = n1803_o[3];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n1822_o = n1820_o | n1821_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n1823_o = n1803_o[2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n1824_o = n1822_o | n1823_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n1825_o = n1803_o[1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n1826_o = n1824_o | n1825_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n1827_o = n1803_o[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n1828_o = n1826_o | n1827_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:223:68  */
  assign n1829_o = ~n1828_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:223:37  */
  assign n1831_o = 1'b1 & n1829_o;
  assign n1836_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:226:9  */
  assign n1837_o = wb_ack_i ? 1'b0 : n1836_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:226:9  */
  assign n1838_o = wb_ack_i ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:223:9  */
  assign n1839_o = n1831_o ? 1'b0 : n1837_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:223:9  */
  assign n1840_o = n1831_o ? 1'b0 : n1838_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:223:9  */
  assign n1841_o = n1831_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:220:9  */
  assign n1842_o = wb_err_i ? 1'b0 : n1839_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:220:9  */
  assign n1843_o = wb_err_i ? 1'b0 : n1840_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:220:9  */
  assign n1844_o = wb_err_i ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:220:9  */
  assign n1845_o = wb_err_i ? 1'b0 : n1841_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:232:59  */
  assign n1846_o = ctrl[114:106];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:232:68  */
  assign n1848_o = n1846_o - 9'b000000001;
  assign n1849_o = {n1848_o, n1845_o, n1844_o, n1843_o};
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:204:7  */
  assign n1850_o = n1786_o ? n1793_o : n1842_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:204:7  */
  assign n1852_o = n1786_o & n1788_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:204:7  */
  assign n1853_o = n1786_o ? 32'b00000000000000000000000000000000 : wb_dat_i;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:204:7  */
  assign n1855_o = n1786_o & n1788_o;
  assign n1856_o = {9'b011111111, 1'b0, 1'b0, 1'b0};
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:204:7  */
  assign n1857_o = n1786_o ? n1856_o : n1849_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:204:7  */
  assign n1859_o = n1786_o & n1788_o;
  assign n1860_o = {n1799_o, n1857_o, n1797_o, n1853_o, n1795_o, n1778_o, n1850_o};
  assign n1862_o = {1'b0, 1'b0, 9'b000000000, 1'b0, 1'b0, 1'b0, 4'b0000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 1'b0, 1'b0, 1'b0};
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:239:17  */
  assign n1865_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2575:36  */
  assign n1872_o = data_i[31:24];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2576:36  */
  assign n1875_o = data_i[23:16];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2577:36  */
  assign n1877_o = data_i[15:8];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2578:36  */
  assign n1879_o = data_i[7:0];
  assign n1880_o = {n1879_o, n1877_o, n1875_o, n1872_o};
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:242:35  */
  assign n1882_o = 1'b0 ? n1880_o : data_i;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2546:42  */
  assign n1889_o = ben_i[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2546:42  */
  assign n1892_o = ben_i[1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2546:42  */
  assign n1894_o = ben_i[2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2546:42  */
  assign n1896_o = ben_i[3];
  assign n1897_o = {n1889_o, n1892_o, n1894_o, n1896_o};
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:243:35  */
  assign n1899_o = 1'b0 ? n1897_o : ben_i;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:247:38  */
  assign n1900_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:247:27  */
  assign n1901_o = n1900_o ? wb_ack_i : 1'b0;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:248:38  */
  assign n1903_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:248:27  */
  assign n1904_o = n1903_o ? wb_dat_i : 32'b00000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:249:23  */
  assign n1906_o = ctrl[98:67];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:249:28  */
  assign n1908_o = 1'b1 ? n1906_o : rdata_gated;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:251:19  */
  assign n1910_o = 1'b1 ? rdata : n1925_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2575:36  */
  assign n1917_o = rdata[31:24];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2576:36  */
  assign n1920_o = rdata[23:16];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2577:36  */
  assign n1922_o = rdata[15:8];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2578:36  */
  assign n1924_o = rdata[7:0];
  assign n1925_o = {n1924_o, n1922_o, n1920_o, n1917_o};
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:252:18  */
  assign n1926_o = ctrl[103];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:252:22  */
  assign n1928_o = 1'b1 ? n1926_o : ack_gated;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:253:18  */
  assign n1929_o = ctrl[104];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:254:18  */
  assign n1930_o = ctrl[105];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:258:25  */
  assign n1932_o = 1'b0 ? priv_i : n1933_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:258:58  */
  assign n1933_o = ctrl[116];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:260:24  */
  assign n1936_o = 1'b0 ? src_i : n1937_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:260:57  */
  assign n1937_o = ctrl[115];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:262:40  */
  assign n1938_o = wren_i | rden_i;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:262:28  */
  assign n1939_o = xbus_access & n1938_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:262:67  */
  assign n1941_o = 1'b0 ? n1939_o : n1945_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:262:101  */
  assign n1942_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:262:121  */
  assign n1943_o = ctrl[1];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:262:112  */
  assign n1944_o = ~n1943_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:262:107  */
  assign n1945_o = n1942_o & n1944_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:263:40  */
  assign n1946_o = wren_i | rden_i;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:263:28  */
  assign n1947_o = xbus_access & n1946_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:263:60  */
  assign n1948_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:263:52  */
  assign n1949_o = n1947_o | n1948_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:263:67  */
  assign n1951_o = 1'b0 ? n1949_o : n1952_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:263:101  */
  assign n1952_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:265:22  */
  assign n1954_o = 1'b0 ? addr_i : n1955_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:265:55  */
  assign n1955_o = ctrl[34:3];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:266:22  */
  assign n1957_o = 1'b0 ? data_i : n1958_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:266:55  */
  assign n1958_o = ctrl[66:35];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:267:32  */
  assign n1959_o = ctrl[2];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:267:44  */
  assign n1960_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:267:35  */
  assign n1961_o = n1959_o & n1960_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:267:23  */
  assign n1962_o = wren_i | n1961_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:267:52  */
  assign n1964_o = 1'b0 ? n1962_o : n1965_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:267:85  */
  assign n1965_o = ctrl[2];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:268:26  */
  assign n1967_o = 1'b0 ? end_byteen : n1968_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:268:59  */
  assign n1968_o = ctrl[102:99];
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:269:23  */
  assign n1970_o = 1'b0 ? stb_int : cyc_int;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:194:5  */
  always @(posedge clk_i or posedge n1763_o)
    if (n1763_o)
      n1971_q <= n1862_o;
    else
      n1971_q <= n1860_o;
  /* ../neorv32/rtl/core/neorv32_wishbone.vhd:180:5  */
  assign n1972_o = {n1936_o, 1'b0, n1932_o};
endmodule

module neorv32_boot_rom_8aaa057a3ce108fd664b4f820549d0c7a5c85d77
  (input  clk_i,
   input  rden_i,
   input  wren_i,
   input  [31:0] addr_i,
   output [31:0] data_o,
   output ack_o,
   output err_o);
  wire acc_en;
  wire rden;
  wire [31:0] rdata;
  wire [9:0] addr;
  wire [16:0] n1677_o;
  wire n1679_o;
  wire n1680_o;
  wire [9:0] n1682_o;
  wire n1685_o;
  wire n1686_o;
  wire [9:0] n1689_o;
  wire [31:0] n1698_o;
  reg n1700_q;
  reg n1703_q;
  reg [31:0] n1705_data; // mem_rd
  assign data_o = n1698_o;
  assign ack_o = rden;
  assign err_o = n1703_q;
  /* ../neorv32/rtl/core/neorv32_boot_rom.vhd:69:10  */
  assign acc_en = n1680_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_boot_rom.vhd:70:10  */
  assign rden = n1700_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_boot_rom.vhd:71:10  */
  assign rdata = n1705_data; // (signal)
  /* ../neorv32/rtl/core/neorv32_boot_rom.vhd:72:10  */
  assign addr = n1682_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_boot_rom.vhd:90:29  */
  assign n1677_o = addr_i[31:15];
  /* ../neorv32/rtl/core/neorv32_boot_rom.vhd:90:56  */
  assign n1679_o = n1677_o == 17'b11111111111111110;
  /* ../neorv32/rtl/core/neorv32_boot_rom.vhd:90:17  */
  assign n1680_o = n1679_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_boot_rom.vhd:91:19  */
  assign n1682_o = addr_i[11:2];
  /* ../neorv32/rtl/core/neorv32_boot_rom.vhd:99:23  */
  assign n1685_o = acc_en & rden_i;
  /* ../neorv32/rtl/core/neorv32_boot_rom.vhd:100:23  */
  assign n1686_o = acc_en & wren_i;
  /* ../neorv32/rtl/core/neorv32_boot_rom.vhd:102:26  */
  assign n1689_o = 10'b1111111111 - addr;
  /* ../neorv32/rtl/core/neorv32_boot_rom.vhd:108:19  */
  assign n1698_o = rden ? rdata : 32'b00000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_boot_rom.vhd:98:5  */
  always @(posedge clk_i)
    n1700_q <= n1685_o;
  /* ../neorv32/rtl/core/neorv32_boot_rom.vhd:98:5  */
  always @(posedge clk_i)
    n1703_q <= n1686_o;
  /* ../neorv32/rtl/core/neorv32_boot_rom.vhd:54:5  */
  reg [31:0] n1704[1023:0] ; // memory
  initial begin
    n1704[1023] = 32'b00110000000000000101000001110011;
    n1704[1022] = 32'b00110000010000000001000001110011;
    n1704[1021] = 32'b00000000000000000000000010010111;
    n1704[1020] = 32'b00001110000000001000000010010011;
    n1704[1019] = 32'b00110000010100001001000001110011;
    n1704[1018] = 32'b10000000000000010000000100010111;
    n1704[1017] = 32'b00011110100000010000000100010011;
    n1704[1016] = 32'b10000000000000010000000110010111;
    n1704[1015] = 32'b01111110010000011000000110010011;
    n1704[1014] = 32'b00000000000000000000001000010011;
    n1704[1013] = 32'b00000000000000000000001010010011;
    n1704[1012] = 32'b00000000000000000000001100010011;
    n1704[1011] = 32'b00000000000000000000001110010011;
    n1704[1010] = 32'b00000000000000000000010000010011;
    n1704[1009] = 32'b00000000000000000000010010010011;
    n1704[1008] = 32'b00000000000000000000100000010011;
    n1704[1007] = 32'b00000000000000000000100010010011;
    n1704[1006] = 32'b00000000000000000000100100010011;
    n1704[1005] = 32'b00000000000000000000100110010011;
    n1704[1004] = 32'b00000000000000000000101000010011;
    n1704[1003] = 32'b00000000000000000000101010010011;
    n1704[1002] = 32'b00000000000000000000101100010011;
    n1704[1001] = 32'b00000000000000000000101110010011;
    n1704[1000] = 32'b00000000000000000000110000010011;
    n1704[999] = 32'b00000000000000000000110010010011;
    n1704[998] = 32'b00000000000000000000110100010011;
    n1704[997] = 32'b00000000000000000000110110010011;
    n1704[996] = 32'b00000000000000000000111000010011;
    n1704[995] = 32'b00000000000000000000111010010011;
    n1704[994] = 32'b00000000000000000000111100010011;
    n1704[993] = 32'b00000000000000000000111110010011;
    n1704[992] = 32'b00000000000000000001010110010111;
    n1704[991] = 32'b11110101000001011000010110010011;
    n1704[990] = 32'b10000000000000010000011000010111;
    n1704[989] = 32'b11110111110001100000011000010011;
    n1704[988] = 32'b10000000000000010000011010010111;
    n1704[987] = 32'b11110111010001101000011010010011;
    n1704[986] = 32'b00000000110001011000111001100011;
    n1704[985] = 32'b00000000110101100101110001100011;
    n1704[984] = 32'b00000000000001011010011100000011;
    n1704[983] = 32'b00000000111001100010000000100011;
    n1704[982] = 32'b00000000010001011000010110010011;
    n1704[981] = 32'b00000000010001100000011000010011;
    n1704[980] = 32'b11111110110111111111000001101111;
    n1704[979] = 32'b10000000000000010000011100010111;
    n1704[978] = 32'b11110101000001110000011100010011;
    n1704[977] = 32'b10000000100000011000011110010011;
    n1704[976] = 32'b00000000111101110101100001100011;
    n1704[975] = 32'b00000000000001110010000000100011;
    n1704[974] = 32'b00000000010001110000011100010011;
    n1704[973] = 32'b11111111010111111111000001101111;
    n1704[972] = 32'b00000000000000000000010100010011;
    n1704[971] = 32'b00000000000000000000010110010011;
    n1704[970] = 32'b00000110000000000000000011101111;
    n1704[969] = 32'b00110000010000000001000001110011;
    n1704[968] = 32'b00110100000001010001000001110011;
    n1704[967] = 32'b00010000010100000000000001110011;
    n1704[966] = 32'b00000000000000000000000001101111;
    n1704[965] = 32'b11111111100000010000000100010011;
    n1704[964] = 32'b00000000100000010010000000100011;
    n1704[963] = 32'b00000000100100010010001000100011;
    n1704[962] = 32'b00110100001000000010010001110011;
    n1704[961] = 32'b00000010000001000100011001100011;
    n1704[960] = 32'b00110100000100000010010001110011;
    n1704[959] = 32'b00000000000001000001010010000011;
    n1704[958] = 32'b00000000001101001111010010010011;
    n1704[957] = 32'b00000000001001000000010000010011;
    n1704[956] = 32'b00110100000101000001000001110011;
    n1704[955] = 32'b00000000001100000000010000010011;
    n1704[954] = 32'b00000000100101000001100001100011;
    n1704[953] = 32'b00110100000100000010010001110011;
    n1704[952] = 32'b00000000001001000000010000010011;
    n1704[951] = 32'b00110100000101000001000001110011;
    n1704[950] = 32'b00000000000000010010010000000011;
    n1704[949] = 32'b00000000010000010010010010000011;
    n1704[948] = 32'b00000000100000010000000100010011;
    n1704[947] = 32'b00110000001000000000000001110011;
    n1704[946] = 32'b11111011000000010000000100010011;
    n1704[945] = 32'b00000100100100010010001000100011;
    n1704[944] = 32'b10000000000000000000010010110111;
    n1704[943] = 32'b00000000000001001010001000100011;
    n1704[942] = 32'b10000000000000000000011110110111;
    n1704[941] = 32'b00000000000001111010000000100011;
    n1704[940] = 32'b11111111111111110001011110110111;
    n1704[939] = 32'b00000100000100010010011000100011;
    n1704[938] = 32'b00000100100000010010010000100011;
    n1704[937] = 32'b00000101001000010010000000100011;
    n1704[936] = 32'b00000011001100010010111000100011;
    n1704[935] = 32'b00000011010000010010110000100011;
    n1704[934] = 32'b00000011010100010010101000100011;
    n1704[933] = 32'b00000011011000010010100000100011;
    n1704[932] = 32'b00000011011100010010011000100011;
    n1704[931] = 32'b00000011100000010010010000100011;
    n1704[930] = 32'b00000011100100010010001000100011;
    n1704[929] = 32'b00000011101000010010000000100011;
    n1704[928] = 32'b00000001101100010010111000100011;
    n1704[927] = 32'b10100011010001111000011110010011;
    n1704[926] = 32'b00110000010101111001000001110011;
    n1704[925] = 32'b11111110100000000010011110000011;
    n1704[924] = 32'b00000000000010000000011100110111;
    n1704[923] = 32'b00000000111001111111011110110011;
    n1704[922] = 32'b00000000000001111000100001100011;
    n1704[921] = 32'b11111010000000000010010000100011;
    n1704[920] = 32'b00010000000100000000011110010011;
    n1704[919] = 32'b11111010111100000010010000100011;
    n1704[918] = 32'b11111110100000000010011110000011;
    n1704[917] = 32'b01000000000000000000011100110111;
    n1704[916] = 32'b00000000111001111111011110110011;
    n1704[915] = 32'b00000110000001111000100001100011;
    n1704[914] = 32'b11110100000000000010000000100011;
    n1704[913] = 32'b11110100000000000010010000100011;
    n1704[912] = 32'b00000000000000000110011110110111;
    n1704[911] = 32'b11110100000000000010011000100011;
    n1704[910] = 32'b00100000010101111000011110010011;
    n1704[909] = 32'b11110100111100000010000000100011;
    n1704[908] = 32'b11110100000000000010010000100011;
    n1704[907] = 32'b11110100000000000010011000100011;
    n1704[906] = 32'b11110100000000000010011110000011;
    n1704[905] = 32'b00000000111001111111011110110011;
    n1704[904] = 32'b11111110000001111001110011100011;
    n1704[903] = 32'b11110100000000000010011110000011;
    n1704[902] = 32'b00000010000000000000011100110111;
    n1704[901] = 32'b00000000111001111110011110110011;
    n1704[900] = 32'b11110100111100000010000000100011;
    n1704[899] = 32'b11110100000000000010011110000011;
    n1704[898] = 32'b00001000000000000000011100110111;
    n1704[897] = 32'b00000000111001111110011110110011;
    n1704[896] = 32'b11110100111100000010000000100011;
    n1704[895] = 32'b11110100000000000010011110000011;
    n1704[894] = 32'b11111110000111111110011100110111;
    n1704[893] = 32'b01000011111101110000011100010011;
    n1704[892] = 32'b00000000111001111111011110110011;
    n1704[891] = 32'b00000000100000000001011100110111;
    n1704[890] = 32'b01100000000001110000011100010011;
    n1704[889] = 32'b00000000111001111110011110110011;
    n1704[888] = 32'b11110100111100000010000000100011;
    n1704[887] = 32'b11111110100000000010011110000011;
    n1704[886] = 32'b00000000000000010000011100110111;
    n1704[885] = 32'b00000000111001111111011110110011;
    n1704[884] = 32'b00000000000001111000100001100011;
    n1704[883] = 32'b00000000000100000000011110010011;
    n1704[882] = 32'b11111100111100000010010000100011;
    n1704[881] = 32'b11111100000000000010011000100011;
    n1704[880] = 32'b11111010000000000010000000100011;
    n1704[879] = 32'b11111110000000000010011010000011;
    n1704[878] = 32'b00000000000000001001011100110111;
    n1704[877] = 32'b11111111111111110111011000110111;
    n1704[876] = 32'b00000000000000000000011110010011;
    n1704[875] = 32'b01011111111101110000011100010011;
    n1704[874] = 32'b10100000000001100000011000010011;
    n1704[873] = 32'b00100000110101110110001001100011;
    n1704[872] = 32'b00000000000000000000011100010011;
    n1704[871] = 32'b00111111111000000000011000010011;
    n1704[870] = 32'b00100000111101100110001001100011;
    n1704[869] = 32'b11111111111101111000011110010011;
    n1704[868] = 32'b00000000000000010000011010110111;
    n1704[867] = 32'b00000000011001111001011110010011;
    n1704[866] = 32'b11111111111101101000011010010011;
    n1704[865] = 32'b00000000001101110001011100010011;
    n1704[864] = 32'b00000001100001110111011100010011;
    n1704[863] = 32'b00000000110101111111011110110011;
    n1704[862] = 32'b00000000111001111110011110110011;
    n1704[861] = 32'b00000000000101111110011110010011;
    n1704[860] = 32'b11111010111100000010000000100011;
    n1704[859] = 32'b11111110100000000010011110000011;
    n1704[858] = 32'b00000000000000100000011100110111;
    n1704[857] = 32'b00000000111001111111011110110011;
    n1704[856] = 32'b00000010000001111000011001100011;
    n1704[855] = 32'b11111000000000000010100000100011;
    n1704[854] = 32'b11111000000000000010101000100011;
    n1704[853] = 32'b11111110000000000010011110000011;
    n1704[852] = 32'b00000000001001111101011110010011;
    n1704[851] = 32'b11111000111100000010110000100011;
    n1704[850] = 32'b11111000000000000010111000100011;
    n1704[849] = 32'b00001000000000000000011110010011;
    n1704[848] = 32'b00110000010001111001000001110011;
    n1704[847] = 32'b00000000100000000000011110010011;
    n1704[846] = 32'b00110000000001111010000001110011;
    n1704[845] = 32'b11111111111111110001010100110111;
    n1704[844] = 32'b11011100010001010000010100010011;
    n1704[843] = 32'b01101011000000000000000011101111;
    n1704[842] = 32'b11110001001100000010010101110011;
    n1704[841] = 32'b01100011010000000000000011101111;
    n1704[840] = 32'b11111111111111110001010100110111;
    n1704[839] = 32'b11011111110001010000010100010011;
    n1704[838] = 32'b01101001110000000000000011101111;
    n1704[837] = 32'b11111110010000000010010100000011;
    n1704[836] = 32'b01100010000000000000000011101111;
    n1704[835] = 32'b11111111111111110001010100110111;
    n1704[834] = 32'b11100000010001010000010100010011;
    n1704[833] = 32'b01101000100000000000000011101111;
    n1704[832] = 32'b11111110000000000010010100000011;
    n1704[831] = 32'b01100000110000000000000011101111;
    n1704[830] = 32'b11111111111111110001010100110111;
    n1704[829] = 32'b11100000110001010000010100010011;
    n1704[828] = 32'b01100111010000000000000011101111;
    n1704[827] = 32'b00110000000100000010010101110011;
    n1704[826] = 32'b01011111100000000000000011101111;
    n1704[825] = 32'b11111111111111110001010100110111;
    n1704[824] = 32'b11100001010001010000010100010011;
    n1704[823] = 32'b01100110000000000000000011101111;
    n1704[822] = 32'b11111100000000000010010101110011;
    n1704[821] = 32'b01011110010000000000000011101111;
    n1704[820] = 32'b11111111111111110001010100110111;
    n1704[819] = 32'b11100001110001010000010100010011;
    n1704[818] = 32'b01100100110000000000000011101111;
    n1704[817] = 32'b11111110100000000010010100000011;
    n1704[816] = 32'b11111111111111110001010000110111;
    n1704[815] = 32'b11111111111111110001100100110111;
    n1704[814] = 32'b01011100100000000000000011101111;
    n1704[813] = 32'b11111111111111110001010100110111;
    n1704[812] = 32'b11100010010001010000010100010011;
    n1704[811] = 32'b01100011000000000000000011101111;
    n1704[810] = 32'b11111111100000000010010100000011;
    n1704[809] = 32'b01011011010000000000000011101111;
    n1704[808] = 32'b11100010110001000000010100010011;
    n1704[807] = 32'b01100010000000000000000011101111;
    n1704[806] = 32'b11111111000000000010010100000011;
    n1704[805] = 32'b01011010010000000000000011101111;
    n1704[804] = 32'b11111111111111110001010100110111;
    n1704[803] = 32'b11100011100001010000010100010011;
    n1704[802] = 32'b01100000110000000000000011101111;
    n1704[801] = 32'b11111111110000000010010100000011;
    n1704[800] = 32'b01011001000000000000000011101111;
    n1704[799] = 32'b11100010110001000000010100010011;
    n1704[798] = 32'b01011111110000000000000011101111;
    n1704[797] = 32'b11111111010000000010010100000011;
    n1704[796] = 32'b01011000000000000000000011101111;
    n1704[795] = 32'b11011100000010010000010100010011;
    n1704[794] = 32'b01011110110000000000000011101111;
    n1704[793] = 32'b11111110100000000010011110000011;
    n1704[792] = 32'b00000000000000100000011100110111;
    n1704[791] = 32'b00000000111001111111011110110011;
    n1704[790] = 32'b00000100000001111000110001100011;
    n1704[789] = 32'b11111111111111110001010100110111;
    n1704[788] = 32'b11100100000001010000010100010011;
    n1704[787] = 32'b01011101000000000000000011101111;
    n1704[786] = 32'b00101011110000000000000011101111;
    n1704[785] = 32'b11111110000000000010010000000011;
    n1704[784] = 32'b00000000000001000000101000110111;
    n1704[783] = 32'b00000000000000010000101010110111;
    n1704[782] = 32'b00000000001101000001010000010011;
    n1704[781] = 32'b00000000101001000000100110110011;
    n1704[780] = 32'b00000000100010011011010000110011;
    n1704[779] = 32'b00000000101101000000010000110011;
    n1704[778] = 32'b11111110100000000010011110000011;
    n1704[777] = 32'b00000001010001111111011110110011;
    n1704[776] = 32'b00001010000001111000011001100011;
    n1704[775] = 32'b11111010000000000010011110000011;
    n1704[774] = 32'b00000001010101111111011110110011;
    n1704[773] = 32'b00001010000001111000000001100011;
    n1704[772] = 32'b11111111111111110001010100110111;
    n1704[771] = 32'b11111010010000000010011110000011;
    n1704[770] = 32'b11100110110001010000010100010011;
    n1704[769] = 32'b01011000100000000000000011101111;
    n1704[768] = 32'b11111111111111110001101000110111;
    n1704[767] = 32'b11100111100010100000010100010011;
    n1704[766] = 32'b01010111110000000000000011101111;
    n1704[765] = 32'b00000110110000000000101010010011;
    n1704[764] = 32'b00000111100000000000101110010011;
    n1704[763] = 32'b00000111001100000000110000010011;
    n1704[762] = 32'b00000110010100000000110010010011;
    n1704[761] = 32'b11111111111111110001011110110111;
    n1704[760] = 32'b11101111100001111000010100010011;
    n1704[759] = 32'b01010110000000000000000011101111;
    n1704[758] = 32'b11111010000000000010011110000011;
    n1704[757] = 32'b00000000000000010000011100110111;
    n1704[756] = 32'b00000000111001111111011110110011;
    n1704[755] = 32'b11111110000001111000101011100011;
    n1704[754] = 32'b11111010010000000010010000000011;
    n1704[753] = 32'b00001111111101000111010000010011;
    n1704[752] = 32'b00000000000001000000010100010011;
    n1704[751] = 32'b01001011010000000000000011101111;
    n1704[750] = 32'b11011100000010010000010100010011;
    n1704[749] = 32'b01010011100000000000000011101111;
    n1704[748] = 32'b00000111001000000000011110010011;
    n1704[747] = 32'b00000110111101000001000001100011;
    n1704[746] = 32'b11111111111111110000001010110111;
    n1704[745] = 32'b00000000000000101000000001100111;
    n1704[744] = 32'b00000000110001101000011010110011;
    n1704[743] = 32'b00000000000101111000011110010011;
    n1704[742] = 32'b11011111010111111111000001101111;
    n1704[741] = 32'b11111111111001110000011010010011;
    n1704[740] = 32'b11111111110101101111011010010011;
    n1704[739] = 32'b00000000000001101001100001100011;
    n1704[738] = 32'b00000000001101111101011110010011;
    n1704[737] = 32'b00000000000101110000011100010011;
    n1704[736] = 32'b11011110100111111111000001101111;
    n1704[735] = 32'b00000000000101111101011110010011;
    n1704[734] = 32'b11111111010111111111000001101111;
    n1704[733] = 32'b00011110100000000000000011101111;
    n1704[732] = 32'b11110100100001011110010011100011;
    n1704[731] = 32'b00000000101101000001010001100011;
    n1704[730] = 32'b11110101001101010110000011100011;
    n1704[729] = 32'b00000000000100000000010100010011;
    n1704[728] = 32'b01110001100000000000000011101111;
    n1704[727] = 32'b11011100000010010000010100010011;
    n1704[726] = 32'b01001101110000000000000011101111;
    n1704[725] = 32'b00000000000000000000010100010011;
    n1704[724] = 32'b00000110100100000000000011101111;
    n1704[723] = 32'b00011001010101000000100001100011;
    n1704[722] = 32'b00000010100010101110010001100011;
    n1704[721] = 32'b00011001100101000000100001100011;
    n1704[720] = 32'b00000110100000000000011110010011;
    n1704[719] = 32'b11100111100010100000010100010011;
    n1704[718] = 32'b00000010111101000000110001100011;
    n1704[717] = 32'b00000011111100000000011110010011;
    n1704[716] = 32'b00011000111101000000110001100011;
    n1704[715] = 32'b11111111111111110001010100110111;
    n1704[714] = 32'b11111001110001010000010100010011;
    n1704[713] = 32'b00000010010000000000000001101111;
    n1704[712] = 32'b00000111010100000000011110010011;
    n1704[711] = 32'b00000010111101000000001001100011;
    n1704[710] = 32'b00010111011101000000110001100011;
    n1704[709] = 32'b11111111100001000001010011100011;
    n1704[708] = 32'b00000000010001001010010000000011;
    n1704[707] = 32'b00000010000001000001000001100011;
    n1704[706] = 32'b11111111111111110001010100110111;
    n1704[705] = 32'b11110000000001010000010100010011;
    n1704[704] = 32'b01001000010000000000000011101111;
    n1704[703] = 32'b11110001100111111111000001101111;
    n1704[702] = 32'b00000000000000000000010100010011;
    n1704[701] = 32'b01101010110000000000000011101111;
    n1704[700] = 32'b11110000110111111111000001101111;
    n1704[699] = 32'b11111111111111110001010100110111;
    n1704[698] = 32'b11110001110001010000010100010011;
    n1704[697] = 32'b01000110100000000000000011101111;
    n1704[696] = 32'b00000000000001000000010100010011;
    n1704[695] = 32'b00111110110000000000000011101111;
    n1704[694] = 32'b11111111111111110001010100110111;
    n1704[693] = 32'b11110010010001010000010100010011;
    n1704[692] = 32'b01000101010000000000000011101111;
    n1704[691] = 32'b00000000010000000000010100110111;
    n1704[690] = 32'b00111101100000000000000011101111;
    n1704[689] = 32'b11111111111111110001010100110111;
    n1704[688] = 32'b11110011110001010000010100010011;
    n1704[687] = 32'b01000100000000000000000011101111;
    n1704[686] = 32'b00000000000000010000011100110111;
    n1704[685] = 32'b11111010000000000010011110000011;
    n1704[684] = 32'b00000000111001111111011110110011;
    n1704[683] = 32'b11111110000001111000110011100011;
    n1704[682] = 32'b11111010010000000010100110000011;
    n1704[681] = 32'b00001111111110011111100110010011;
    n1704[680] = 32'b00000000000010011000010100010011;
    n1704[679] = 32'b00111001010000000000000011101111;
    n1704[678] = 32'b00000111100100000000011110010011;
    n1704[677] = 32'b11101010111110011001100011100011;
    n1704[676] = 32'b00101010000000000000000011101111;
    n1704[675] = 32'b00000000000001010000011001100011;
    n1704[674] = 32'b00000000001100000000010100010011;
    n1704[673] = 32'b01000110000000000000000011101111;
    n1704[672] = 32'b11111111111111110001010100110111;
    n1704[671] = 32'b11110100100001010000010100010011;
    n1704[670] = 32'b00111111110000000000000011101111;
    n1704[669] = 32'b00000001000001000101101100010011;
    n1704[668] = 32'b00000000010000000000100110110111;
    n1704[667] = 32'b00000000000000010000110110110111;
    n1704[666] = 32'b11111111111100000000110100010011;
    n1704[665] = 32'b00100010000000000000000011101111;
    n1704[664] = 32'b00010101000000000000000011101111;
    n1704[663] = 32'b00001101100000000000010100010011;
    n1704[662] = 32'b00001111010000000000000011101111;
    n1704[661] = 32'b00000000000010011000010100010011;
    n1704[660] = 32'b00010000010000000000000011101111;
    n1704[659] = 32'b00001101010000000000000011101111;
    n1704[658] = 32'b00100010010000000000000011101111;
    n1704[657] = 32'b00000000000101010111010100010011;
    n1704[656] = 32'b11111110000001010001110011100011;
    n1704[655] = 32'b11111111111110110000101100010011;
    n1704[654] = 32'b00000001101110011000100110110011;
    n1704[653] = 32'b11111101101010110001100011100011;
    n1704[652] = 32'b11111111000000000010011010000011;
    n1704[651] = 32'b00000000010000000000100110110111;
    n1704[650] = 32'b00000000000000000000110100010011;
    n1704[649] = 32'b00000000000000000000110110010011;
    n1704[648] = 32'b00000000110010011000011110010011;
    n1704[647] = 32'b00000000110111010000011100110011;
    n1704[646] = 32'b00000000000001110010010110000011;
    n1704[645] = 32'b00000000111111010000010100110011;
    n1704[644] = 32'b00000000110100010010011000100011;
    n1704[643] = 32'b00000000101111011000110110110011;
    n1704[642] = 32'b00100110110000000000000011101111;
    n1704[641] = 32'b00000000010000000000011110110111;
    n1704[640] = 32'b00000000010011010000110100010011;
    n1704[639] = 32'b00000000110000010010011010000011;
    n1704[638] = 32'b00000000110001111000011110010011;
    n1704[637] = 32'b11111100100011010110110011100011;
    n1704[636] = 32'b01000111100010001101010110110111;
    n1704[635] = 32'b10101111111001011000010110010011;
    n1704[634] = 32'b00000000010000000000010100110111;
    n1704[633] = 32'b00100100100000000000000011101111;
    n1704[632] = 32'b00000000000001000000010110010011;
    n1704[631] = 32'b00000000010010011000010100010011;
    n1704[630] = 32'b00100011110000000000000011101111;
    n1704[629] = 32'b00000000100010011000010100010011;
    n1704[628] = 32'b01000001101100000000010110110011;
    n1704[627] = 32'b00100011000000000000000011101111;
    n1704[626] = 32'b11111111111111110001010100110111;
    n1704[625] = 32'b11011010100001010000010100010011;
    n1704[624] = 32'b11101100000111111111000001101111;
    n1704[623] = 32'b00000000000100000000010100010011;
    n1704[622] = 32'b11101100010111111111000001101111;
    n1704[621] = 32'b00000000010001001010011110000011;
    n1704[620] = 32'b11100100000001111001111011100011;
    n1704[619] = 32'b11111111111111110001010100110111;
    n1704[618] = 32'b11110101100001010000010100010011;
    n1704[617] = 32'b11101010010111111111000001101111;
    n1704[616] = 32'b00000000000100000000010100010011;
    n1704[615] = 32'b11100100110111111111000001101111;
    n1704[614] = 32'b11111111111111110001010100110111;
    n1704[613] = 32'b11110110100001010000010100010011;
    n1704[612] = 32'b11101001000111111111000001101111;
    n1704[611] = 32'b11111001010000000010010110000011;
    n1704[610] = 32'b11111001000000000010010100000011;
    n1704[609] = 32'b11111001010000000010011110000011;
    n1704[608] = 32'b11111110111101011001101011100011;
    n1704[607] = 32'b00000000000000001000000001100111;
    n1704[606] = 32'b11111010100000000000011100010011;
    n1704[605] = 32'b00000000000001110010011110000011;
    n1704[604] = 32'b11111011111101111111011110010011;
    n1704[603] = 32'b00000000111101110010000000100011;
    n1704[602] = 32'b00000000000000001000000001100111;
    n1704[601] = 32'b11111010101000000010011000100011;
    n1704[600] = 32'b11111010100000000010011110000011;
    n1704[599] = 32'b11111110000001111100111011100011;
    n1704[598] = 32'b11111010110000000010010100000011;
    n1704[597] = 32'b00001111111101010111010100010011;
    n1704[596] = 32'b00000000000000001000000001100111;
    n1704[595] = 32'b11111111000000010000000100010011;
    n1704[594] = 32'b00000000100000010010010000100011;
    n1704[593] = 32'b00000000000001010000010000010011;
    n1704[592] = 32'b00000001000001010101010100010011;
    n1704[591] = 32'b00001111111101010111010100010011;
    n1704[590] = 32'b00000000000100010010011000100011;
    n1704[589] = 32'b11111101000111111111000011101111;
    n1704[588] = 32'b00000000100001000101010100010011;
    n1704[587] = 32'b00001111111101010111010100010011;
    n1704[586] = 32'b11111100010111111111000011101111;
    n1704[585] = 32'b00001111111101000111010100010011;
    n1704[584] = 32'b00000000100000010010010000000011;
    n1704[583] = 32'b00000000110000010010000010000011;
    n1704[582] = 32'b00000001000000010000000100010011;
    n1704[581] = 32'b11111011000111111111000001101111;
    n1704[580] = 32'b11111010100000000000011100010011;
    n1704[579] = 32'b00000000000001110010011110000011;
    n1704[578] = 32'b11111000011101111111011110010011;
    n1704[577] = 32'b00000100000001111110011110010011;
    n1704[576] = 32'b00000000111101110010000000100011;
    n1704[575] = 32'b00000000000000001000000001100111;
    n1704[574] = 32'b11111101000000010000000100010011;
    n1704[573] = 32'b00000010100100010010001000100011;
    n1704[572] = 32'b00000011001000010010000000100011;
    n1704[571] = 32'b00000001001100010010111000100011;
    n1704[570] = 32'b00000001010000010010110000100011;
    n1704[569] = 32'b00000001010100010010101000100011;
    n1704[568] = 32'b00000010000100010010011000100011;
    n1704[567] = 32'b00000010100000010010010000100011;
    n1704[566] = 32'b00000000000001010000100100010011;
    n1704[565] = 32'b00000000000001011000100110010011;
    n1704[564] = 32'b00000000000000000000010010010011;
    n1704[563] = 32'b00000000000000010000101010110111;
    n1704[562] = 32'b00000000010000000000101000010011;
    n1704[561] = 32'b00000100000010010001101001100011;
    n1704[560] = 32'b11111010000000000010011110000011;
    n1704[559] = 32'b00000001010101111111011110110011;
    n1704[558] = 32'b11111110000001111000110011100011;
    n1704[557] = 32'b11111010010000000010010000000011;
    n1704[556] = 32'b00001111111101000111010000010011;
    n1704[555] = 32'b00000000110000010000011110010011;
    n1704[554] = 32'b00000000100101111000011110110011;
    n1704[553] = 32'b00000000100001111000000000100011;
    n1704[552] = 32'b00000000000101001000010010010011;
    n1704[551] = 32'b11111101010001001001110011100011;
    n1704[550] = 32'b00000010110000010010000010000011;
    n1704[549] = 32'b00000010100000010010010000000011;
    n1704[548] = 32'b00000000110000010010010100000011;
    n1704[547] = 32'b00000010010000010010010010000011;
    n1704[546] = 32'b00000010000000010010100100000011;
    n1704[545] = 32'b00000001110000010010100110000011;
    n1704[544] = 32'b00000001100000010010101000000011;
    n1704[543] = 32'b00000001010000010010101010000011;
    n1704[542] = 32'b00000011000000010000000100010011;
    n1704[541] = 32'b00000000000000001000000001100111;
    n1704[540] = 32'b11110110000111111111000011101111;
    n1704[539] = 32'b00000000001100000000010100010011;
    n1704[538] = 32'b00000000100110011000010000110011;
    n1704[537] = 32'b11110000000111111111000011101111;
    n1704[536] = 32'b00000000000001000000010100010011;
    n1704[535] = 32'b11110001000111111111000011101111;
    n1704[534] = 32'b00000000000000000000010100010011;
    n1704[533] = 32'b11101111000111111111000011101111;
    n1704[532] = 32'b00000000000001010000010000010011;
    n1704[531] = 32'b11101101010111111111000011101111;
    n1704[530] = 32'b11111001110111111111000001101111;
    n1704[529] = 32'b11111111000000010000000100010011;
    n1704[528] = 32'b00000000000100010010011000100011;
    n1704[527] = 32'b11110010110111111111000011101111;
    n1704[526] = 32'b00000000011000000000010100010011;
    n1704[525] = 32'b11101101000111111111000011101111;
    n1704[524] = 32'b00000000110000010010000010000011;
    n1704[523] = 32'b00000001000000010000000100010011;
    n1704[522] = 32'b11101011000111111111000001101111;
    n1704[521] = 32'b11111110000000010000000100010011;
    n1704[520] = 32'b00000000000100010010111000100011;
    n1704[519] = 32'b11110000110111111111000011101111;
    n1704[518] = 32'b00000000010100000000010100010011;
    n1704[517] = 32'b11101011000111111111000011101111;
    n1704[516] = 32'b00000000000000000000010100010011;
    n1704[515] = 32'b11101010100111111111000011101111;
    n1704[514] = 32'b00000000101000010010011000100011;
    n1704[513] = 32'b11101000110111111111000011101111;
    n1704[512] = 32'b00000001110000010010000010000011;
    n1704[511] = 32'b00000000110000010010010100000011;
    n1704[510] = 32'b00000010000000010000000100010011;
    n1704[509] = 32'b00000000000000001000000001100111;
    n1704[508] = 32'b11111111000000010000000100010011;
    n1704[507] = 32'b00000000000100010010011000100011;
    n1704[506] = 32'b11101101100111111111000011101111;
    n1704[505] = 32'b00001010101100000000010100010011;
    n1704[504] = 32'b11100111110111111111000011101111;
    n1704[503] = 32'b11100110010111111111000011101111;
    n1704[502] = 32'b11111001010111111111000011101111;
    n1704[501] = 32'b11111011000111111111000011101111;
    n1704[500] = 32'b00000000001001010111011110010011;
    n1704[499] = 32'b11111111111100000000010100010011;
    n1704[498] = 32'b00000010000001111000000001100011;
    n1704[497] = 32'b11101011010111111111000011101111;
    n1704[496] = 32'b00000000010000000000010100010011;
    n1704[495] = 32'b11100101100111111111000011101111;
    n1704[494] = 32'b11100100000111111111000011101111;
    n1704[493] = 32'b11111001000111111111000011101111;
    n1704[492] = 32'b00000001111001010001010100010011;
    n1704[491] = 32'b01000001111101010101010100010011;
    n1704[490] = 32'b00000000110000010010000010000011;
    n1704[489] = 32'b00000001000000010000000100010011;
    n1704[488] = 32'b00000000000000001000000001100111;
    n1704[487] = 32'b11111101000000010000000100010011;
    n1704[486] = 32'b00000010100000010010010000100011;
    n1704[485] = 32'b00000010100100010010001000100011;
    n1704[484] = 32'b00000001001100010010111000100011;
    n1704[483] = 32'b00000010000100010010011000100011;
    n1704[482] = 32'b00000011001000010010000000100011;
    n1704[481] = 32'b00000001010000010010110000100011;
    n1704[480] = 32'b00000000000001010000010010010011;
    n1704[479] = 32'b00000000101100010010011000100011;
    n1704[478] = 32'b00000000000000000000010000010011;
    n1704[477] = 32'b00000000010000000000100110010011;
    n1704[476] = 32'b00000000110000010000011110010011;
    n1704[475] = 32'b00000000100001111000011110110011;
    n1704[474] = 32'b00000000000001111100101000000011;
    n1704[473] = 32'b11110010000111111111000011101111;
    n1704[472] = 32'b11100101000111111111000011101111;
    n1704[471] = 32'b00000000001000000000010100010011;
    n1704[470] = 32'b11011111010111111111000011101111;
    n1704[469] = 32'b00000000100001001000100100110011;
    n1704[468] = 32'b00000000000010010000010100010011;
    n1704[467] = 32'b11100000000111111111000011101111;
    n1704[466] = 32'b00000000000010100000010100010011;
    n1704[465] = 32'b11011110000111111111000011101111;
    n1704[464] = 32'b11011100100111111111000011101111;
    n1704[463] = 32'b11110001100111111111000011101111;
    n1704[462] = 32'b00000000000101010111010100010011;
    n1704[461] = 32'b11111110000001010001110011100011;
    n1704[460] = 32'b00000000000101000000010000010011;
    n1704[459] = 32'b11111011001101000001111011100011;
    n1704[458] = 32'b00000010110000010010000010000011;
    n1704[457] = 32'b00000010100000010010010000000011;
    n1704[456] = 32'b00000010010000010010010010000011;
    n1704[455] = 32'b00000010000000010010100100000011;
    n1704[454] = 32'b00000001110000010010100110000011;
    n1704[453] = 32'b00000001100000010010101000000011;
    n1704[452] = 32'b00000011000000010000000100010011;
    n1704[451] = 32'b00000000000000001000000001100111;
    n1704[450] = 32'b00000000001000000000011100110111;
    n1704[449] = 32'b11111010000000000010011110000011;
    n1704[448] = 32'b00000000111001111111011110110011;
    n1704[447] = 32'b11111110000001111001110011100011;
    n1704[446] = 32'b11111010101000000010001000100011;
    n1704[445] = 32'b00000000000000001000000001100111;
    n1704[444] = 32'b11111110000000010000000100010011;
    n1704[443] = 32'b00000001001000010010100000100011;
    n1704[442] = 32'b00000000000001010000100100010011;
    n1704[441] = 32'b00000011000000000000010100010011;
    n1704[440] = 32'b00000000000100010010111000100011;
    n1704[439] = 32'b00000000100000010010110000100011;
    n1704[438] = 32'b00000000100100010010101000100011;
    n1704[437] = 32'b00000001001100010010011000100011;
    n1704[436] = 32'b11111100100111111111000011101111;
    n1704[435] = 32'b00000111100000000000010100010011;
    n1704[434] = 32'b11111111111111110001010010110111;
    n1704[433] = 32'b11111011110111111111000011101111;
    n1704[432] = 32'b00000001110000000000010000010011;
    n1704[431] = 32'b11111010100001001000010010010011;
    n1704[430] = 32'b11111111110000000000100110010011;
    n1704[429] = 32'b00000000100010010101011110110011;
    n1704[428] = 32'b00000000111101111111011110010011;
    n1704[427] = 32'b00000000111101001000011110110011;
    n1704[426] = 32'b00000000000001111100010100000011;
    n1704[425] = 32'b11111111110001000000010000010011;
    n1704[424] = 32'b11111001100111111111000011101111;
    n1704[423] = 32'b11111111001101000001010011100011;
    n1704[422] = 32'b00000001110000010010000010000011;
    n1704[421] = 32'b00000001100000010010010000000011;
    n1704[420] = 32'b00000001010000010010010010000011;
    n1704[419] = 32'b00000001000000010010100100000011;
    n1704[418] = 32'b00000000110000010010100110000011;
    n1704[417] = 32'b00000010000000010000000100010011;
    n1704[416] = 32'b00000000000000001000000001100111;
    n1704[415] = 32'b11111111000000010000000100010011;
    n1704[414] = 32'b00000000100000010010010000100011;
    n1704[413] = 32'b00000001001000010010000000100011;
    n1704[412] = 32'b00000000000100010010011000100011;
    n1704[411] = 32'b00000000100100010010001000100011;
    n1704[410] = 32'b00000000000001010000010000010011;
    n1704[409] = 32'b00000000101000000000100100010011;
    n1704[408] = 32'b00000000000001000100010010000011;
    n1704[407] = 32'b00000000000101000000010000010011;
    n1704[406] = 32'b00000000000001001001111001100011;
    n1704[405] = 32'b00000000110000010010000010000011;
    n1704[404] = 32'b00000000100000010010010000000011;
    n1704[403] = 32'b00000000010000010010010010000011;
    n1704[402] = 32'b00000000000000010010100100000011;
    n1704[401] = 32'b00000001000000010000000100010011;
    n1704[400] = 32'b00000000000000001000000001100111;
    n1704[399] = 32'b00000001001001001001011001100011;
    n1704[398] = 32'b00000000110100000000010100010011;
    n1704[397] = 32'b11110010110111111111000011101111;
    n1704[396] = 32'b00000000000001001000010100010011;
    n1704[395] = 32'b11110010010111111111000011101111;
    n1704[394] = 32'b11111100100111111111000001101111;
    n1704[393] = 32'b11111111000000010000000100010011;
    n1704[392] = 32'b00000000100000010010010000100011;
    n1704[391] = 32'b00000000000001010000010000010011;
    n1704[390] = 32'b11111111111111110001010100110111;
    n1704[389] = 32'b11010110000001010000010100010011;
    n1704[388] = 32'b00000000000100010010011000100011;
    n1704[387] = 32'b11111001000111111111000011101111;
    n1704[386] = 32'b00000000001001000001011110010011;
    n1704[385] = 32'b11111111111111110001010100110111;
    n1704[384] = 32'b00000000100001111000011110110011;
    n1704[383] = 32'b11111011100001010000010100010011;
    n1704[382] = 32'b00000000111101010000010100110011;
    n1704[381] = 32'b11110111100111111111000011101111;
    n1704[380] = 32'b00000000100000000000011110010011;
    n1704[379] = 32'b00110000000001111011000001110011;
    n1704[378] = 32'b11111110100000000010011110000011;
    n1704[377] = 32'b00000000000000010000011100110111;
    n1704[376] = 32'b00000000111001111111011110110011;
    n1704[375] = 32'b00000000000001111000100001100011;
    n1704[374] = 32'b00000000000100000000011110010011;
    n1704[373] = 32'b11111100111100000010010000100011;
    n1704[372] = 32'b11111100000000000010011000100011;
    n1704[371] = 32'b00000000000000000000000001101111;
    n1704[370] = 32'b11111011000000010000000100010011;
    n1704[369] = 32'b00000100000100010010011000100011;
    n1704[368] = 32'b00000100010100010010010000100011;
    n1704[367] = 32'b00000100011000010010001000100011;
    n1704[366] = 32'b00000100011100010010000000100011;
    n1704[365] = 32'b00000010100000010010111000100011;
    n1704[364] = 32'b00000010100100010010110000100011;
    n1704[363] = 32'b00000010101000010010101000100011;
    n1704[362] = 32'b00000010101100010010100000100011;
    n1704[361] = 32'b00000010110000010010011000100011;
    n1704[360] = 32'b00000010110100010010010000100011;
    n1704[359] = 32'b00000010111000010010001000100011;
    n1704[358] = 32'b00000010111100010010000000100011;
    n1704[357] = 32'b00000001000000010010111000100011;
    n1704[356] = 32'b00000001000100010010110000100011;
    n1704[355] = 32'b00000001110000010010101000100011;
    n1704[354] = 32'b00000001110100010010100000100011;
    n1704[353] = 32'b00000001111000010010011000100011;
    n1704[352] = 32'b00000001111100010010010000100011;
    n1704[351] = 32'b00110100001000000010010011110011;
    n1704[350] = 32'b10000000000000000000011110110111;
    n1704[349] = 32'b00000000011101111000011110010011;
    n1704[348] = 32'b00001010111101001001011001100011;
    n1704[347] = 32'b11111110100000000010011110000011;
    n1704[346] = 32'b00000000000000010000011100110111;
    n1704[345] = 32'b00000000111001111111011110110011;
    n1704[344] = 32'b00000000000001111000100001100011;
    n1704[343] = 32'b11111100100000000010011110000011;
    n1704[342] = 32'b00000000000101111100011110010011;
    n1704[341] = 32'b11111100111100000010010000100011;
    n1704[340] = 32'b11111110100000000010011110000011;
    n1704[339] = 32'b00000000000000100000011100110111;
    n1704[338] = 32'b00000000111001111111011110110011;
    n1704[337] = 32'b00000010000001111000100001100011;
    n1704[336] = 32'b10111011010111111111000011101111;
    n1704[335] = 32'b11111110000000000010011110000011;
    n1704[334] = 32'b11111111111100000000011100010011;
    n1704[333] = 32'b11111000111000000010110000100011;
    n1704[332] = 32'b00000000001001111101011110010011;
    n1704[331] = 32'b00000000101001111000010100110011;
    n1704[330] = 32'b00000000111101010011011110110011;
    n1704[329] = 32'b00000000101101111000011110110011;
    n1704[328] = 32'b11111000111100000010111000100011;
    n1704[327] = 32'b11111000101000000010110000100011;
    n1704[326] = 32'b00000000000000000000000000010011;
    n1704[325] = 32'b00000011110000010010010000000011;
    n1704[324] = 32'b00000100110000010010000010000011;
    n1704[323] = 32'b00000100100000010010001010000011;
    n1704[322] = 32'b00000100010000010010001100000011;
    n1704[321] = 32'b00000100000000010010001110000011;
    n1704[320] = 32'b00000011100000010010010010000011;
    n1704[319] = 32'b00000011010000010010010100000011;
    n1704[318] = 32'b00000011000000010010010110000011;
    n1704[317] = 32'b00000010110000010010011000000011;
    n1704[316] = 32'b00000010100000010010011010000011;
    n1704[315] = 32'b00000010010000010010011100000011;
    n1704[314] = 32'b00000010000000010010011110000011;
    n1704[313] = 32'b00000001110000010010100000000011;
    n1704[312] = 32'b00000001100000010010100010000011;
    n1704[311] = 32'b00000001010000010010111000000011;
    n1704[310] = 32'b00000001000000010010111010000011;
    n1704[309] = 32'b00000000110000010010111100000011;
    n1704[308] = 32'b00000000100000010010111110000011;
    n1704[307] = 32'b00000101000000010000000100010011;
    n1704[306] = 32'b00110000001000000000000001110011;
    n1704[305] = 32'b00000000011100000000011110010011;
    n1704[304] = 32'b00000000111101001001110001100011;
    n1704[303] = 32'b10000000000000000000011110110111;
    n1704[302] = 32'b00000000000001111010011110000011;
    n1704[301] = 32'b00000000000001111000011001100011;
    n1704[300] = 32'b00000000000100000000010100010011;
    n1704[299] = 32'b11101000100111111111000011101111;
    n1704[298] = 32'b00110100000100000010010001110011;
    n1704[297] = 32'b11111110100000000010011110000011;
    n1704[296] = 32'b00000000000001000000011100110111;
    n1704[295] = 32'b00000000111001111111011110110011;
    n1704[294] = 32'b00000100000001111000001001100011;
    n1704[293] = 32'b11111111111111110001010100110111;
    n1704[292] = 32'b11010110100001010000010100010011;
    n1704[291] = 32'b11100001000111111111000011101111;
    n1704[290] = 32'b00000000000001001000010100010011;
    n1704[289] = 32'b11011001010111111111000011101111;
    n1704[288] = 32'b00000010000000000000010100010011;
    n1704[287] = 32'b11010111010111111111000011101111;
    n1704[286] = 32'b00000000000001000000010100010011;
    n1704[285] = 32'b11011000010111111111000011101111;
    n1704[284] = 32'b00000010000000000000010100010011;
    n1704[283] = 32'b11010110010111111111000011101111;
    n1704[282] = 32'b00110100001100000010010101110011;
    n1704[281] = 32'b11010111010111111111000011101111;
    n1704[280] = 32'b11111111111111110001010100110111;
    n1704[279] = 32'b11011100000001010000010100010011;
    n1704[278] = 32'b11011101110111111111000011101111;
    n1704[277] = 32'b00000000010001000000010000010011;
    n1704[276] = 32'b00110100000101000001000001110011;
    n1704[275] = 32'b11110011100111111111000001101111;
    n1704[274] = 32'b11111101000000010000000100010011;
    n1704[273] = 32'b00000001011000010010100000100011;
    n1704[272] = 32'b00000000000100000000011110010011;
    n1704[271] = 32'b10000000000000000000101100110111;
    n1704[270] = 32'b00000010100000010010010000100011;
    n1704[269] = 32'b00000010000100010010011000100011;
    n1704[268] = 32'b00000010100100010010001000100011;
    n1704[267] = 32'b00000011001000010010000000100011;
    n1704[266] = 32'b00000001001100010010111000100011;
    n1704[265] = 32'b00000001010000010010110000100011;
    n1704[264] = 32'b00000001010100010010101000100011;
    n1704[263] = 32'b00000001011100010010011000100011;
    n1704[262] = 32'b00000001100000010010010000100011;
    n1704[261] = 32'b00000000111110110010000000100011;
    n1704[260] = 32'b00000000000001010000010000010011;
    n1704[259] = 32'b00000010000001010001100001100011;
    n1704[258] = 32'b11111111111111110001010100110111;
    n1704[257] = 32'b11010111010001010000010100010011;
    n1704[256] = 32'b11011000010111111111000011101111;
    n1704[255] = 32'b00000000010000000000010110110111;
    n1704[254] = 32'b00000000000001000000010100010011;
    n1704[253] = 32'b10101111110111111111000011101111;
    n1704[252] = 32'b01000111100010001101011110110111;
    n1704[251] = 32'b10101111111001111000011110010011;
    n1704[250] = 32'b00000100111101010000100001100011;
    n1704[249] = 32'b00000000000000000000010100010011;
    n1704[248] = 32'b00000011100000000000000001101111;
    n1704[247] = 32'b11111111111111110001010100110111;
    n1704[246] = 32'b11011001010001010000010100010011;
    n1704[245] = 32'b11010101100111111111000011101111;
    n1704[244] = 32'b00000000010000000000010100110111;
    n1704[243] = 32'b11001101110111111111000011101111;
    n1704[242] = 32'b11111111111111110001010100110111;
    n1704[241] = 32'b11011010000001010000010100010011;
    n1704[240] = 32'b11010100010111111111000011101111;
    n1704[239] = 32'b11111110100000000010011110000011;
    n1704[238] = 32'b00000000000010000000011100110111;
    n1704[237] = 32'b00000000111001111111011110110011;
    n1704[236] = 32'b00000000000001111001011001100011;
    n1704[235] = 32'b00000000001100000000010100010011;
    n1704[234] = 32'b11011000010111111111000011101111;
    n1704[233] = 32'b10111011010111111111000011101111;
    n1704[232] = 32'b11111010000001010000001011100011;
    n1704[231] = 32'b11111111000111111111000001101111;
    n1704[230] = 32'b00000000010000000000100110110111;
    n1704[229] = 32'b00000000010010011000010110010011;
    n1704[228] = 32'b00000000000001000000010100010011;
    n1704[227] = 32'b10101001010111111111000011101111;
    n1704[226] = 32'b00000000000001010000101000010011;
    n1704[225] = 32'b00000000100010011000010110010011;
    n1704[224] = 32'b00000000000001000000010100010011;
    n1704[223] = 32'b10101000010111111111000011101111;
    n1704[222] = 32'b11111111000000000010110000000011;
    n1704[221] = 32'b00000000000001010000101010010011;
    n1704[220] = 32'b11111111110010100111101110010011;
    n1704[219] = 32'b00000000000000000000100100010011;
    n1704[218] = 32'b00000000000000000000010010010011;
    n1704[217] = 32'b00000000110010011000100110010011;
    n1704[216] = 32'b00000001001110010000010110110011;
    n1704[215] = 32'b00000101011110010001110001100011;
    n1704[214] = 32'b00000001010101001000010010110011;
    n1704[213] = 32'b00000000001000000000010100010011;
    n1704[212] = 32'b11111010000001001001010011100011;
    n1704[211] = 32'b11111111111111110001010100110111;
    n1704[210] = 32'b11011010100001010000010100010011;
    n1704[209] = 32'b11001100100111111111000011101111;
    n1704[208] = 32'b00000010110000010010000010000011;
    n1704[207] = 32'b00000010100000010010010000000011;
    n1704[206] = 32'b10000000000000000000011110110111;
    n1704[205] = 32'b00000001010001111010001000100011;
    n1704[204] = 32'b00000000000010110010000000100011;
    n1704[203] = 32'b00000010010000010010010010000011;
    n1704[202] = 32'b00000010000000010010100100000011;
    n1704[201] = 32'b00000001110000010010100110000011;
    n1704[200] = 32'b00000001100000010010101000000011;
    n1704[199] = 32'b00000001010000010010101010000011;
    n1704[198] = 32'b00000001000000010010101100000011;
    n1704[197] = 32'b00000000110000010010101110000011;
    n1704[196] = 32'b00000000100000010010110000000011;
    n1704[195] = 32'b00000011000000010000000100010011;
    n1704[194] = 32'b00000000000000001000000001100111;
    n1704[193] = 32'b00000000000001000000010100010011;
    n1704[192] = 32'b10100000100111111111000011101111;
    n1704[191] = 32'b00000001001011000000011110110011;
    n1704[190] = 32'b00000000101001001000010010110011;
    n1704[189] = 32'b00000000101001111010000000100011;
    n1704[188] = 32'b00000000010010010000100100010011;
    n1704[187] = 32'b11111000110111111111000001101111;
    n1704[186] = 32'b11111111000000010000000100010011;
    n1704[185] = 32'b00000000000100010010011000100011;
    n1704[184] = 32'b00000000100000010010010000100011;
    n1704[183] = 32'b00000000100000000000011110010011;
    n1704[182] = 32'b00110000000001111011000001110011;
    n1704[181] = 32'b11111111000000000010010000000011;
    n1704[180] = 32'b00000000000001010000010001100011;
    n1704[179] = 32'b01000000010000000000010000110111;
    n1704[178] = 32'b11111111111111110001010100110111;
    n1704[177] = 32'b11011010110001010000010100010011;
    n1704[176] = 32'b11000100010111111111000011101111;
    n1704[175] = 32'b00000000000001000000010100010011;
    n1704[174] = 32'b10111100100111111111000011101111;
    n1704[173] = 32'b11111111111111110001010100110111;
    n1704[172] = 32'b11011011110001010000010100010011;
    n1704[171] = 32'b11000011000111111111000011101111;
    n1704[170] = 32'b11111010000000000010011110000011;
    n1704[169] = 32'b11111110000001111100111011100011;
    n1704[168] = 32'b00000000000001000000000011100111;
    n1704[167] = 32'b01010010010001010000101000000111;
    n1704[166] = 32'b00000000000000000101111101010010;
    n1704[165] = 32'b01010010010100100100010100001010;
    n1704[164] = 32'b01000011010110000100010101011111;
    n1704[163] = 32'b00000000000000000000000000100000;
    n1704[162] = 32'b01101001011000010111011101000001;
    n1704[161] = 32'b01100111011011100110100101110100;
    n1704[160] = 32'b01101111011001010110111000100000;
    n1704[159] = 32'b00110010001100110111011001110010;
    n1704[158] = 32'b01100101011110000110010101011111;
    n1704[157] = 32'b01101110011010010110001000101110;
    n1704[156] = 32'b00100000001011100010111000101110;
    n1704[155] = 32'b00000000000000000000000000000000;
    n1704[154] = 32'b01100100011000010110111101001100;
    n1704[153] = 32'b00100000011001110110111001101001;
    n1704[152] = 32'b00000000000000000100000000101000;
    n1704[151] = 32'b00101110001011100010111000101001;
    n1704[150] = 32'b00000000000000000000000000001010;
    n1704[149] = 32'b00000000000000000100101101001111;
    n1704[148] = 32'b01110100011011110110111101000010;
    n1704[147] = 32'b00100000011001110110111001101001;
    n1704[146] = 32'b01101101011011110111001001100110;
    n1704[145] = 32'b00000000000000000000000000100000;
    n1704[144] = 32'b00001010001011100010111000101110;
    n1704[143] = 32'b00000000000000000000000000001010;
    n1704[142] = 32'b00111100000010100000101000001010;
    n1704[141] = 32'b01000101010011100010000000111100;
    n1704[140] = 32'b00110011010101100101001001001111;
    n1704[139] = 32'b01101111010000100010000000110010;
    n1704[138] = 32'b01101111011011000111010001101111;
    n1704[137] = 32'b01110010011001010110010001100001;
    n1704[136] = 32'b00001010001111100011111000100000;
    n1704[135] = 32'b01000100010011000100001000001010;
    n1704[134] = 32'b01001101001000000011101001010110;
    n1704[133] = 32'b00110001001000000111001001100001;
    n1704[132] = 32'b00110000001100100010000000110110;
    n1704[131] = 32'b01001000000010100011001100110010;
    n1704[130] = 32'b00100000001110100101011001010111;
    n1704[129] = 32'b00000000000000000000000000100000;
    n1704[128] = 32'b01000100010010010100001100001010;
    n1704[127] = 32'b00000000001000000010000000111010;
    n1704[126] = 32'b01001011010011000100001100001010;
    n1704[125] = 32'b00000000001000000010000000111010;
    n1704[124] = 32'b01010011010010010100110100001010;
    n1704[123] = 32'b00000000001000000011101001000001;
    n1704[122] = 32'b01010011010010010101100000001010;
    n1704[121] = 32'b00000000001000000011101001000001;
    n1704[120] = 32'b01000011010011110101001100001010;
    n1704[119] = 32'b00000000001000000010000000111010;
    n1704[118] = 32'b01000101010011010100100100001010;
    n1704[117] = 32'b00000000001000000011101001001101;
    n1704[116] = 32'b01110100011110010110001000100000;
    n1704[115] = 32'b01000000001000000111001101100101;
    n1704[114] = 32'b00000000000000000000000000000000;
    n1704[113] = 32'b01000101010011010100010000001010;
    n1704[112] = 32'b00000000001000000011101001001101;
    n1704[111] = 32'b01110100011101010100000100001010;
    n1704[110] = 32'b01101111011011110110001001101111;
    n1704[109] = 32'b01101110011010010010000001110100;
    n1704[108] = 32'b00101110011100110011100000100000;
    n1704[107] = 32'b01100101011100100101000000100000;
    n1704[106] = 32'b01100001001000000111001101110011;
    n1704[105] = 32'b01101011001000000111100101101110;
    n1704[104] = 32'b01110100001000000111100101100101;
    n1704[103] = 32'b01100010011000010010000001101111;
    n1704[102] = 32'b00101110011101000111001001101111;
    n1704[101] = 32'b00000000000000000000000000001010;
    n1704[100] = 32'b01110010011011110110001001000001;
    n1704[99] = 32'b00101110011001000110010101110100;
    n1704[98] = 32'b00000000000000000000101000001010;
    n1704[97] = 32'b01101001011000010111011001000001;
    n1704[96] = 32'b01101100011000100110000101101100;
    n1704[95] = 32'b01001101010000110010000001100101;
    n1704[94] = 32'b00001010001110100111001101000100;
    n1704[93] = 32'b00100000001110100110100000100000;
    n1704[92] = 32'b01110000011011000110010101001000;
    n1704[91] = 32'b00111010011100100010000000001010;
    n1704[90] = 32'b01110011011001010101001000100000;
    n1704[89] = 32'b01110100011100100110000101110100;
    n1704[88] = 32'b00111010011101010010000000001010;
    n1704[87] = 32'b01101100011100000101010100100000;
    n1704[86] = 32'b00001010011001000110000101101111;
    n1704[85] = 32'b00100000001110100111001100100000;
    n1704[84] = 32'b01110010011011110111010001010011;
    n1704[83] = 32'b01101111011101000010000001100101;
    n1704[82] = 32'b01100001011011000110011000100000;
    n1704[81] = 32'b00100000000010100110100001110011;
    n1704[80] = 32'b01001100001000000011101001101100;
    n1704[79] = 32'b00100000011001000110000101101111;
    n1704[78] = 32'b01101101011011110111001001100110;
    n1704[77] = 32'b01100001011011000110011000100000;
    n1704[76] = 32'b00100000000010100110100001110011;
    n1704[75] = 32'b01000010001000000011101001111000;
    n1704[74] = 32'b00100000011101000110111101101111;
    n1704[73] = 32'b01101101011011110111001001100110;
    n1704[72] = 32'b01100001011011000110011000100000;
    n1704[71] = 32'b00101000001000000110100001110011;
    n1704[70] = 32'b00101001010100000100100101011000;
    n1704[69] = 32'b00111010011001010010000000001010;
    n1704[68] = 32'b01100101011110000100010100100000;
    n1704[67] = 32'b01100101011101000111010101100011;
    n1704[66] = 32'b00000000000000000000000000000000;
    n1704[65] = 32'b01000100010011010100001100001010;
    n1704[64] = 32'b00000000001000000011111000111010;
    n1704[63] = 32'b01100101001000000110111101001110;
    n1704[62] = 32'b01110101011000110110010101111000;
    n1704[61] = 32'b01101100011000100110000101110100;
    n1704[60] = 32'b01110110011000010010000001100101;
    n1704[59] = 32'b01100001011011000110100101100001;
    n1704[58] = 32'b00101110011001010110110001100010;
    n1704[57] = 32'b00000000000000000000000000000000;
    n1704[56] = 32'b01110100011010010111001001010111;
    n1704[55] = 32'b00000000000000000010000001100101;
    n1704[54] = 32'b01110100011110010110001000100000;
    n1704[53] = 32'b01110100001000000111001101100101;
    n1704[52] = 32'b01010000010100110010000001101111;
    n1704[51] = 32'b01101100011001100010000001001001;
    n1704[50] = 32'b00100000011010000111001101100001;
    n1704[49] = 32'b00000000000000000010000001000000;
    n1704[48] = 32'b01111001001010000010000000111111;
    n1704[47] = 32'b00100000001010010110111000101111;
    n1704[46] = 32'b00000000000000000000000000000000;
    n1704[45] = 32'b01100001011011000100011000001010;
    n1704[44] = 32'b01101110011010010110100001110011;
    n1704[43] = 32'b00101110001011100010111001100111;
    n1704[42] = 32'b00000000000000000000000000100000;
    n1704[41] = 32'b01100101001000000110111101001110;
    n1704[40] = 32'b01110101011000110110010101111000;
    n1704[39] = 32'b01101100011000100110000101110100;
    n1704[38] = 32'b00000000000000000010111001100101;
    n1704[37] = 32'b00100000001010010110001100101000;
    n1704[36] = 32'b01010011001000000111100101100010;
    n1704[35] = 32'b01101000011100000110010101110100;
    n1704[34] = 32'b01001110001000000110111001100001;
    n1704[33] = 32'b01101001011101000110110001101111;
    n1704[32] = 32'b01100111000010100110011101101110;
    n1704[31] = 32'b01110101011010000111010001101001;
    n1704[30] = 32'b01101111011000110010111001100010;
    n1704[29] = 32'b01110100011100110010111101101101;
    n1704[28] = 32'b01110100011011000110111101101110;
    n1704[27] = 32'b00101111011001110110111001101001;
    n1704[26] = 32'b01110010011011110110010101101110;
    n1704[25] = 32'b00000000001100100011001101110110;
    n1704[24] = 32'b01100001011101100110111001001001;
    n1704[23] = 32'b00100000011001000110100101101100;
    n1704[22] = 32'b00000000010001000100110101000011;
    n1704[21] = 32'b00110011001100100011000100110000;
    n1704[20] = 32'b00110111001101100011010100110100;
    n1704[19] = 32'b01100010011000010011100100111000;
    n1704[18] = 32'b01100110011001010110010001100011;
    n1704[17] = 32'b00000000010001010101100001000101;
    n1704[16] = 32'b01011010010010010101001100000000;
    n1704[15] = 32'b01001000010000110000000001000101;
    n1704[14] = 32'b01000110000000000101001101001011;
    n1704[13] = 32'b00000000010010000101001101001100;
    n1704[12] = 32'b00000000000000000000000000000000;
    n1704[11] = 32'b00000000000000000000000000000000;
    n1704[10] = 32'b00000000000000000000000000000000;
    n1704[9] = 32'b00000000000000000000000000000000;
    n1704[8] = 32'b00000000000000000000000000000000;
    n1704[7] = 32'b00000000000000000000000000000000;
    n1704[6] = 32'b00000000000000000000000000000000;
    n1704[5] = 32'b00000000000000000000000000000000;
    n1704[4] = 32'b00000000000000000000000000000000;
    n1704[3] = 32'b00000000000000000000000000000000;
    n1704[2] = 32'b00000000000000000000000000000000;
    n1704[1] = 32'b00000000000000000000000000000000;
    n1704[0] = 32'b00000000000000000000000000000000;
    end
  always @(posedge clk_i)
    if (acc_en)
      n1705_data <= n1704[n1689_o];
  /* ../neorv32/rtl/core/neorv32_boot_rom.vhd:98:5  */
endmodule

module neorv32_dmem_2048_34d7de1b571aa545cf571b84dc4b40d1f42fed39
  (input  clk_i,
   input  rden_i,
   input  wren_i,
   input  [3:0] ben_i,
   input  [31:0] addr_i,
   input  [31:0] data_i,
   output [31:0] data_o,
   output ack_o);
  wire acc_en;
  wire [31:0] rdata;
  wire rden;
  wire [8:0] addr;
  wire [8:0] addr_ff;
  wire [7:0] mem_ram_b0_rd;
  wire [7:0] mem_ram_b1_rd;
  wire [7:0] mem_ram_b2_rd;
  wire [7:0] mem_ram_b3_rd;
  wire [20:0] n1566_o;
  wire n1568_o;
  wire n1569_o;
  wire [8:0] n1572_o;
  wire n1575_o;
  wire n1576_o;
  wire [7:0] n1581_o;
  wire n1584_o;
  wire n1585_o;
  wire [7:0] n1590_o;
  wire n1593_o;
  wire n1594_o;
  wire [7:0] n1599_o;
  wire n1602_o;
  wire n1603_o;
  wire [7:0] n1608_o;
  wire n1611_o;
  wire n1612_o;
  wire n1613_o;
  wire n1614_o;
  wire n1643_o;
  wire n1644_o;
  wire n1645_o;
  wire [15:0] n1649_o;
  wire [23:0] n1650_o;
  wire [31:0] n1651_o;
  wire [31:0] n1652_o;
  reg n1654_q;
  reg [8:0] n1655_q;
  reg n1664_q;
  wire [7:0] n1665_data; // mem_rd
  wire [7:0] n1667_data; // mem_rd
  wire [7:0] n1669_data; // mem_rd
  wire [7:0] n1671_data; // mem_rd
  assign data_o = n1652_o;
  assign ack_o = n1664_q;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:49:10  */
  assign acc_en = n1569_o; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:50:10  */
  assign rdata = n1651_o; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:51:10  */
  assign rden = n1654_q; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:52:10  */
  assign addr = n1572_o; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:53:10  */
  assign addr_ff = n1655_q; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:67:10  */
  assign mem_ram_b0_rd = n1665_data; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:67:25  */
  assign mem_ram_b1_rd = n1667_data; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:67:40  */
  assign mem_ram_b2_rd = n1669_data; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:67:55  */
  assign mem_ram_b3_rd = n1671_data; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:83:29  */
  assign n1566_o = addr_i[31:11];
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:83:56  */
  assign n1568_o = n1566_o == 21'b100000000000000000000;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:83:17  */
  assign n1569_o = n1568_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:84:19  */
  assign n1572_o = addr_i[10:2];
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:94:37  */
  assign n1575_o = ben_i[0];
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:94:27  */
  assign n1576_o = wren_i & n1575_o;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:95:59  */
  assign n1581_o = data_i[7:0];
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:97:37  */
  assign n1584_o = ben_i[1];
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:97:27  */
  assign n1585_o = wren_i & n1584_o;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:98:59  */
  assign n1590_o = data_i[15:8];
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:100:37  */
  assign n1593_o = ben_i[2];
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:100:27  */
  assign n1594_o = wren_i & n1593_o;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:101:59  */
  assign n1599_o = data_i[23:16];
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:103:37  */
  assign n1602_o = ben_i[3];
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:103:27  */
  assign n1603_o = wren_i & n1602_o;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:104:59  */
  assign n1608_o = data_i[31:24];
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:93:7  */
  assign n1611_o = acc_en & n1576_o;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:93:7  */
  assign n1612_o = acc_en & n1585_o;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:93:7  */
  assign n1613_o = acc_en & n1594_o;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:93:7  */
  assign n1614_o = acc_en & n1603_o;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:122:23  */
  assign n1643_o = acc_en & rden_i;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:123:35  */
  assign n1644_o = rden_i | wren_i;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:123:23  */
  assign n1645_o = acc_en & n1644_o;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:128:26  */
  assign n1649_o = {mem_ram_b3_rd, mem_ram_b2_rd};
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:128:42  */
  assign n1650_o = {n1649_o, mem_ram_b1_rd};
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:128:58  */
  assign n1651_o = {n1650_o, mem_ram_b0_rd};
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:131:19  */
  assign n1652_o = rden ? rdata : 32'b00000000000000000000000000000000;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:121:5  */
  always @(posedge clk_i)
    n1654_q <= n1643_o;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:91:5  */
  always @(posedge clk_i)
    n1655_q <= addr;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:121:5  */
  always @(posedge clk_i)
    n1664_q <= n1645_o;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:111:31  */
  reg [7:0] mem_ram_b0[511:0] ; // memory
  assign n1665_data = mem_ram_b0[addr_ff];
  always @(posedge clk_i)
    if (n1611_o)
      mem_ram_b0[addr] <= n1581_o;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:111:31  */
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:95:22  */
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:112:31  */
  reg [7:0] mem_ram_b1[511:0] ; // memory
  assign n1667_data = mem_ram_b1[addr_ff];
  always @(posedge clk_i)
    if (n1612_o)
      mem_ram_b1[addr] <= n1590_o;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:112:31  */
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:98:22  */
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:113:31  */
  reg [7:0] mem_ram_b2[511:0] ; // memory
  assign n1669_data = mem_ram_b2[addr_ff];
  always @(posedge clk_i)
    if (n1613_o)
      mem_ram_b2[addr] <= n1599_o;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:113:31  */
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:101:22  */
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:114:31  */
  reg [7:0] mem_ram_b3[511:0] ; // memory
  assign n1671_data = mem_ram_b3[addr_ff];
  always @(posedge clk_i)
    if (n1614_o)
      mem_ram_b3[addr] <= n1608_o;
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:114:31  */
  /* ../neorv32/rtl/core/mem/neorv32_dmem.legacy.vhd:104:22  */
endmodule

module neorv32_imem_1024_91a7f356ca6ce41b6122bd41e60c1f2eb8f0f0e3
  (input  clk_i,
   input  rden_i,
   input  wren_i,
   input  [3:0] ben_i,
   input  [31:0] addr_i,
   input  [31:0] data_i,
   output [31:0] data_o,
   output ack_o,
   output err_o);
  wire acc_en;
  wire [31:0] rdata;
  wire rden;
  wire [7:0] addr;
  wire [7:0] addr_ff;
  wire [7:0] mem_b0_rd;
  wire [7:0] mem_b1_rd;
  wire [7:0] mem_b2_rd;
  wire [7:0] mem_b3_rd;
  wire [21:0] n1452_o;
  wire n1454_o;
  wire n1455_o;
  wire [7:0] n1458_o;
  wire n1461_o;
  wire n1462_o;
  wire [7:0] n1467_o;
  wire n1470_o;
  wire n1471_o;
  wire [7:0] n1476_o;
  wire n1479_o;
  wire n1480_o;
  wire [7:0] n1485_o;
  wire n1488_o;
  wire n1489_o;
  wire [7:0] n1494_o;
  wire n1497_o;
  wire n1498_o;
  wire n1499_o;
  wire n1500_o;
  wire [15:0] n1527_o;
  wire [23:0] n1528_o;
  wire [31:0] n1529_o;
  wire n1532_o;
  wire n1533_o;
  wire n1534_o;
  wire [31:0] n1540_o;
  reg n1542_q;
  reg [7:0] n1543_q;
  reg n1553_q;
  reg n1554_q;
  wire [7:0] n1555_data; // mem_rd
  wire [7:0] n1557_data; // mem_rd
  wire [7:0] n1559_data; // mem_rd
  wire [7:0] n1561_data; // mem_rd
  assign data_o = n1540_o;
  assign ack_o = n1553_q;
  assign err_o = n1554_q;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:53:10  */
  assign acc_en = n1455_o; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:54:10  */
  assign rdata = n1529_o; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:55:10  */
  assign rden = n1542_q; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:56:10  */
  assign addr = n1458_o; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:57:10  */
  assign addr_ff = n1543_q; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:84:10  */
  assign mem_b0_rd = n1555_data; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:84:21  */
  assign mem_b1_rd = n1557_data; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:84:32  */
  assign mem_b2_rd = n1559_data; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:84:43  */
  assign mem_b3_rd = n1561_data; // (signal)
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:108:29  */
  assign n1452_o = addr_i[31:10];
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:108:56  */
  assign n1454_o = n1452_o == 22'b0000000000000000000000;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:108:17  */
  assign n1455_o = n1454_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:109:19  */
  assign n1458_o = addr_i[9:2];
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:138:39  */
  assign n1461_o = ben_i[0];
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:138:29  */
  assign n1462_o = wren_i & n1461_o;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:139:61  */
  assign n1467_o = data_i[7:0];
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:141:39  */
  assign n1470_o = ben_i[1];
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:141:29  */
  assign n1471_o = wren_i & n1470_o;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:142:61  */
  assign n1476_o = data_i[15:8];
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:144:39  */
  assign n1479_o = ben_i[2];
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:144:29  */
  assign n1480_o = wren_i & n1479_o;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:145:61  */
  assign n1485_o = data_i[23:16];
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:147:39  */
  assign n1488_o = ben_i[3];
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:147:29  */
  assign n1489_o = wren_i & n1488_o;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:148:61  */
  assign n1494_o = data_i[31:24];
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:137:9  */
  assign n1497_o = acc_en & n1462_o;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:137:9  */
  assign n1498_o = acc_en & n1471_o;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:137:9  */
  assign n1499_o = acc_en & n1480_o;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:137:9  */
  assign n1500_o = acc_en & n1489_o;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:159:24  */
  assign n1527_o = {mem_b3_rd, mem_b2_rd};
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:159:36  */
  assign n1528_o = {n1527_o, mem_b1_rd};
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:159:48  */
  assign n1529_o = {n1528_o, mem_b0_rd};
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:168:22  */
  assign n1532_o = acc_en & rden_i;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:173:37  */
  assign n1533_o = rden_i | wren_i;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:173:25  */
  assign n1534_o = acc_en & n1533_o;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:180:19  */
  assign n1540_o = rden ? rdata : 32'b00000000000000000000000000000000;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:167:5  */
  always @(posedge clk_i)
    n1542_q <= n1532_o;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:135:7  */
  always @(posedge clk_i)
    n1543_q <= addr;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:167:5  */
  always @(posedge clk_i)
    n1553_q <= n1534_o;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:167:5  */
  always @(posedge clk_i)
    n1554_q <= 1'b0;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:154:29  */
  reg [7:0] mem_ram_b0[255:0] ; // memory
  assign n1555_data = mem_ram_b0[addr_ff];
  always @(posedge clk_i)
    if (n1497_o)
      mem_ram_b0[addr] <= n1467_o;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:154:29  */
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:139:24  */
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:155:29  */
  reg [7:0] mem_ram_b1[255:0] ; // memory
  assign n1557_data = mem_ram_b1[addr_ff];
  always @(posedge clk_i)
    if (n1498_o)
      mem_ram_b1[addr] <= n1476_o;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:155:29  */
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:142:24  */
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:156:29  */
  reg [7:0] mem_ram_b2[255:0] ; // memory
  assign n1559_data = mem_ram_b2[addr_ff];
  always @(posedge clk_i)
    if (n1499_o)
      mem_ram_b2[addr] <= n1485_o;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:156:29  */
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:145:24  */
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:157:29  */
  reg [7:0] mem_ram_b3[255:0] ; // memory
  assign n1561_data = mem_ram_b3[addr_ff];
  always @(posedge clk_i)
    if (n1500_o)
      mem_ram_b3[addr] <= n1494_o;
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:157:29  */
  /* ../neorv32/rtl/core/mem/neorv32_imem.legacy.vhd:148:24  */
endmodule

module neorv32_bus_keeper
  (input  clk_i,
   input  rstn_i,
   input  [31:0] addr_i,
   input  rden_i,
   input  wren_i,
   input  [31:0] data_i,
   input  [31:0] bus_addr_i,
   input  bus_rden_i,
   input  bus_wren_i,
   input  bus_ack_i,
   input  bus_err_i,
   input  bus_tmo_i,
   input  bus_ext_i,
   input  bus_xip_i,
   output [31:0] data_o,
   output ack_o,
   output err_o);
  wire err_flag;
  wire err_type;
  wire acc_en;
  wire wren;
  wire rden;
  wire [8:0] control;
  wire [5:0] n1311_o;
  wire n1313_o;
  wire n1314_o;
  wire n1316_o;
  wire n1317_o;
  wire n1319_o;
  wire n1321_o;
  wire n1322_o;
  wire n1323_o;
  wire n1325_o;
  wire n1327_o;
  wire n1338_o;
  wire n1340_o;
  wire n1342_o;
  localparam [31:0] n1343_o = 32'b00000000000000000000000000000000;
  wire [29:0] n1345_o;
  wire [31:0] n1346_o;
  wire n1351_o;
  wire n1359_o;
  wire n1360_o;
  wire n1363_o;
  wire n1365_o;
  wire n1366_o;
  wire n1367_o;
  wire n1368_o;
  wire [3:0] n1369_o;
  wire [3:0] n1371_o;
  wire [3:0] n1372_o;
  wire [3:0] n1373_o;
  wire n1374_o;
  wire n1375_o;
  wire n1376_o;
  wire n1380_o;
  wire n1381_o;
  wire n1382_o;
  wire n1383_o;
  wire n1384_o;
  wire [1:0] n1391_o;
  wire n1392_o;
  wire n1393_o;
  wire n1394_o;
  wire [1:0] n1395_o;
  wire [1:0] n1396_o;
  wire [1:0] n1397_o;
  wire n1398_o;
  wire [1:0] n1399_o;
  wire [1:0] n1400_o;
  wire n1401_o;
  wire [1:0] n1402_o;
  wire [7:0] n1403_o;
  wire [4:0] n1404_o;
  wire [4:0] n1405_o;
  wire [4:0] n1406_o;
  wire [1:0] n1407_o;
  wire n1408_o;
  wire [1:0] n1409_o;
  wire [1:0] n1410_o;
  wire n1411_o;
  wire n1412_o;
  wire [7:0] n1413_o;
  wire [7:0] n1416_o;
  wire [3:0] n1421_o;
  wire n1427_o;
  wire n1429_o;
  wire n1431_o;
  wire n1432_o;
  wire n1433_o;
  wire n1434_o;
  wire n1435_o;
  wire n1436_o;
  wire n1437_o;
  wire n1438_o;
  wire n1440_o;
  reg n1441_q;
  wire n1442_o;
  reg n1443_q;
  reg [7:0] n1444_q;
  wire [8:0] n1445_o;
  reg [31:0] n1446_q;
  reg n1447_q;
  assign data_o = n1446_q;
  assign ack_o = n1447_q;
  assign err_o = n1440_o;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:85:10  */
  assign err_flag = n1441_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:86:10  */
  assign err_type = n1443_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:89:10  */
  assign acc_en = n1314_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:90:10  */
  assign wren = n1316_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:91:10  */
  assign rden = n1317_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:105:10  */
  assign control = n1445_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:119:29  */
  assign n1311_o = addr_i[8:3];
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:119:56  */
  assign n1313_o = n1311_o == 6'b101111;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:119:17  */
  assign n1314_o = n1313_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:120:20  */
  assign n1316_o = acc_en & wren_i;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:121:20  */
  assign n1317_o = acc_en & rden_i;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:126:16  */
  assign n1319_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:130:19  */
  assign n1321_o = control[6];
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:132:29  */
  assign n1322_o = control[5];
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:133:26  */
  assign n1323_o = wren | rden;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:133:7  */
  assign n1325_o = n1323_o ? 1'b0 : err_flag;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:130:7  */
  assign n1327_o = n1321_o ? 1'b1 : n1325_o;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:143:22  */
  assign n1338_o = wren | rden;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:145:7  */
  assign n1340_o = rden ? err_type : 1'b0;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:145:7  */
  assign n1342_o = rden ? err_flag : 1'b0;
  assign n1345_o = n1343_o[30:1];
  assign n1346_o = {n1342_o, n1345_o, n1340_o};
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:157:16  */
  assign n1351_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:168:19  */
  assign n1359_o = control[0];
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:168:27  */
  assign n1360_o = ~n1359_o;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:171:31  */
  assign n1363_o = bus_rden_i | bus_wren_i;
  assign n1365_o = control[0];
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:171:9  */
  assign n1366_o = n1363_o ? 1'b1 : n1365_o;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:177:21  */
  assign n1367_o = control[8];
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:177:29  */
  assign n1368_o = ~n1367_o;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:178:65  */
  assign n1369_o = control[4:1];
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:178:74  */
  assign n1371_o = n1369_o - 4'b0001;
  assign n1372_o = control[4:1];
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:177:9  */
  assign n1373_o = n1368_o ? n1371_o : n1372_o;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:181:35  */
  assign n1374_o = control[7];
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:181:56  */
  assign n1375_o = bus_ext_i | bus_xip_i;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:181:42  */
  assign n1376_o = n1374_o | n1375_o;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:187:25  */
  assign n1380_o = control[8];
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:187:53  */
  assign n1381_o = control[7];
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:187:60  */
  assign n1382_o = ~n1381_o;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:187:40  */
  assign n1383_o = n1380_o & n1382_o;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:187:68  */
  assign n1384_o = n1383_o | bus_tmo_i;
  assign n1391_o = {1'b0, 1'b0};
  assign n1392_o = control[0];
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:192:9  */
  assign n1393_o = bus_ack_i ? 1'b0 : n1392_o;
  assign n1394_o = control[5];
  assign n1395_o = {1'b0, n1394_o};
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:192:9  */
  assign n1396_o = bus_ack_i ? n1391_o : n1395_o;
  assign n1397_o = {1'b1, 1'b1};
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:187:9  */
  assign n1398_o = n1384_o ? 1'b0 : n1393_o;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:187:9  */
  assign n1399_o = n1384_o ? n1397_o : n1396_o;
  assign n1400_o = {1'b1, 1'b0};
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:183:9  */
  assign n1401_o = bus_err_i ? 1'b0 : n1398_o;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:183:9  */
  assign n1402_o = bus_err_i ? n1400_o : n1399_o;
  assign n1403_o = {n1376_o, n1402_o, n1373_o, n1401_o};
  assign n1404_o = {4'b1110, n1366_o};
  assign n1405_o = n1403_o[4:0];
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:168:7  */
  assign n1406_o = n1360_o ? n1404_o : n1405_o;
  assign n1407_o = n1403_o[6:5];
  assign n1408_o = control[5];
  assign n1409_o = {1'b0, n1408_o};
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:168:7  */
  assign n1410_o = n1360_o ? n1409_o : n1407_o;
  assign n1411_o = n1403_o[7];
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:168:7  */
  assign n1412_o = n1360_o ? 1'b0 : n1411_o;
  assign n1413_o = {n1412_o, n1410_o, n1406_o};
  assign n1416_o = {1'b0, 1'b0, 1'b0, 4'b0000, 1'b0};
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:202:52  */
  assign n1421_o = control[4:1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n1427_o = n1421_o[3];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n1429_o = 1'b0 | n1427_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n1431_o = n1421_o[2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n1432_o = n1429_o | n1431_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n1433_o = n1421_o[1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n1434_o = n1432_o | n1433_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n1435_o = n1421_o[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n1436_o = n1434_o | n1435_o;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:202:61  */
  assign n1437_o = ~n1436_o;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:202:26  */
  assign n1438_o = n1437_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:205:20  */
  assign n1440_o = control[6];
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:129:5  */
  always @(posedge clk_i or posedge n1319_o)
    if (n1319_o)
      n1441_q <= 1'b0;
    else
      n1441_q <= n1327_o;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:129:5  */
  assign n1442_o = n1321_o ? n1322_o : err_type;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:129:5  */
  always @(posedge clk_i or posedge n1319_o)
    if (n1319_o)
      n1443_q <= 1'b0;
    else
      n1443_q <= n1442_o;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:163:5  */
  always @(posedge clk_i or posedge n1351_o)
    if (n1351_o)
      n1444_q <= n1416_o;
    else
      n1444_q <= n1413_o;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:157:5  */
  assign n1445_o = {n1438_o, n1444_q};
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:142:5  */
  always @(posedge clk_i)
    n1446_q <= n1346_o;
  /* ../neorv32/rtl/core/neorv32_bus_keeper.vhd:142:5  */
  always @(posedge clk_i)
    n1447_q <= n1338_o;
endmodule

module neorv32_busswitch_3f29546453678b855931c174a97d6c0894b8f546
  (input  clk_i,
   input  rstn_i,
   input  ca_bus_priv_i,
   input  ca_bus_cached_i,
   input  [31:0] ca_bus_addr_i,
   input  [31:0] ca_bus_wdata_i,
   input  [3:0] ca_bus_ben_i,
   input  ca_bus_we_i,
   input  ca_bus_re_i,
   input  cb_bus_priv_i,
   input  cb_bus_cached_i,
   input  [31:0] cb_bus_addr_i,
   input  [31:0] cb_bus_wdata_i,
   input  [3:0] cb_bus_ben_i,
   input  cb_bus_we_i,
   input  cb_bus_re_i,
   input  [31:0] p_bus_rdata_i,
   input  p_bus_ack_i,
   input  p_bus_err_i,
   output [31:0] ca_bus_rdata_o,
   output ca_bus_ack_o,
   output ca_bus_err_o,
   output [31:0] cb_bus_rdata_o,
   output cb_bus_ack_o,
   output cb_bus_err_o,
   output p_bus_priv_o,
   output p_bus_cached_o,
   output p_bus_src_o,
   output [31:0] p_bus_addr_o,
   output [31:0] p_bus_wdata_o,
   output [3:0] p_bus_ben_o,
   output p_bus_we_o,
   output p_bus_re_o);
  wire ca_rd_req_buf;
  wire ca_wr_req_buf;
  wire cb_rd_req_buf;
  wire cb_wr_req_buf;
  wire ca_req_current;
  wire ca_req_pending;
  wire cb_req_current;
  wire cb_req_pending;
  wire ca_bus_ack;
  wire cb_bus_ack;
  wire ca_bus_err;
  wire cb_bus_err;
  wire p_bus_we;
  wire p_bus_re;
  wire [8:0] arbiter;
  wire n1139_o;
  wire [2:0] n1142_o;
  wire n1143_o;
  wire n1144_o;
  wire n1145_o;
  wire n1146_o;
  wire n1147_o;
  wire n1148_o;
  wire n1149_o;
  wire n1150_o;
  wire n1153_o;
  wire n1154_o;
  wire n1155_o;
  wire n1156_o;
  wire n1157_o;
  wire n1158_o;
  wire n1159_o;
  wire n1160_o;
  wire n1161_o;
  wire n1164_o;
  wire n1181_o;
  wire n1183_o;
  wire n1184_o;
  wire n1186_o;
  wire n1187_o;
  wire n1189_o;
  wire n1190_o;
  wire n1192_o;
  wire [2:0] n1194_o;
  wire [2:0] n1198_o;
  wire [3:0] n1207_o;
  wire [3:0] n1208_o;
  wire [3:0] n1209_o;
  wire [3:0] n1210_o;
  wire [3:0] n1211_o;
  wire [3:0] n1212_o;
  wire [3:0] n1213_o;
  wire [3:0] n1214_o;
  wire [3:0] n1215_o;
  wire n1217_o;
  wire n1219_o;
  wire n1220_o;
  wire [2:0] n1223_o;
  wire [2:0] n1224_o;
  wire n1226_o;
  wire n1230_o;
  wire n1232_o;
  wire n1233_o;
  wire [2:0] n1236_o;
  wire [2:0] n1237_o;
  wire n1239_o;
  wire n1243_o;
  wire [4:0] n1245_o;
  wire [2:0] n1246_o;
  reg [2:0] n1247_o;
  wire n1248_o;
  reg n1249_o;
  reg n1250_o;
  reg n1251_o;
  wire n1253_o;
  wire n1254_o;
  wire [31:0] n1255_o;
  wire [31:0] n1257_o;
  wire [31:0] n1259_o;
  wire n1260_o;
  wire n1261_o;
  wire [31:0] n1262_o;
  wire [3:0] n1264_o;
  wire [3:0] n1266_o;
  wire n1267_o;
  wire n1268_o;
  wire [3:0] n1269_o;
  wire n1270_o;
  wire n1271_o;
  wire n1272_o;
  wire n1273_o;
  wire n1274_o;
  wire n1275_o;
  wire n1276_o;
  wire n1277_o;
  wire n1278_o;
  wire n1279_o;
  wire n1280_o;
  wire n1281_o;
  wire n1282_o;
  wire n1283_o;
  wire n1284_o;
  wire n1285_o;
  wire n1286_o;
  wire n1287_o;
  wire n1288_o;
  wire n1289_o;
  wire n1291_o;
  wire n1292_o;
  wire n1294_o;
  wire n1295_o;
  wire n1296_o;
  wire n1298_o;
  wire n1299_o;
  reg n1301_q;
  reg n1302_q;
  reg n1303_q;
  reg n1304_q;
  reg [2:0] n1305_q;
  wire [8:0] n1306_o;
  assign ca_bus_rdata_o = p_bus_rdata_i;
  assign ca_bus_ack_o = ca_bus_ack;
  assign ca_bus_err_o = ca_bus_err;
  assign cb_bus_rdata_o = p_bus_rdata_i;
  assign cb_bus_ack_o = cb_bus_ack;
  assign cb_bus_err_o = cb_bus_err;
  assign p_bus_priv_o = n1275_o;
  assign p_bus_cached_o = n1272_o;
  assign p_bus_src_o = n1286_o;
  assign p_bus_addr_o = n1255_o;
  assign p_bus_wdata_o = n1257_o;
  assign p_bus_ben_o = n1264_o;
  assign p_bus_we_o = n1283_o;
  assign p_bus_re_o = n1285_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:94:10  */
  assign ca_rd_req_buf = n1301_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:94:26  */
  assign ca_wr_req_buf = n1302_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:95:10  */
  assign cb_rd_req_buf = n1303_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:95:26  */
  assign cb_wr_req_buf = n1304_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:96:10  */
  assign ca_req_current = n1183_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:96:26  */
  assign ca_req_pending = n1189_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:97:10  */
  assign cb_req_current = n1186_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:97:26  */
  assign cb_req_pending = n1192_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:100:10  */
  assign ca_bus_ack = n1289_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:100:22  */
  assign cb_bus_ack = n1292_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:101:10  */
  assign ca_bus_err = n1296_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:101:22  */
  assign cb_bus_err = n1299_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:102:10  */
  assign p_bus_we = n1278_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:102:22  */
  assign p_bus_re = n1281_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:113:10  */
  assign arbiter = n1306_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:121:16  */
  assign n1139_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:128:32  */
  assign n1142_o = arbiter[5:3];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:130:39  */
  assign n1143_o = ca_rd_req_buf | ca_bus_re_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:130:76  */
  assign n1144_o = ca_bus_err | ca_bus_ack;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:130:60  */
  assign n1145_o = ~n1144_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:130:55  */
  assign n1146_o = n1143_o & n1145_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:131:39  */
  assign n1147_o = ca_wr_req_buf | ca_bus_we_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:131:76  */
  assign n1148_o = ca_bus_err | ca_bus_ack;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:131:60  */
  assign n1149_o = ~n1148_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:131:55  */
  assign n1150_o = n1147_o & n1149_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:131:92  */
  assign n1153_o = n1150_o & 1'b1;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:133:39  */
  assign n1154_o = cb_rd_req_buf | cb_bus_re_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:133:76  */
  assign n1155_o = cb_bus_err | cb_bus_ack;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:133:60  */
  assign n1156_o = ~n1155_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:133:55  */
  assign n1157_o = n1154_o & n1156_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:134:39  */
  assign n1158_o = cb_wr_req_buf | cb_bus_we_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:134:76  */
  assign n1159_o = cb_bus_err | cb_bus_ack;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:134:60  */
  assign n1160_o = ~n1159_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:134:55  */
  assign n1161_o = n1158_o & n1160_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:134:92  */
  assign n1164_o = n1161_o & 1'b0;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:139:34  */
  assign n1181_o = ca_bus_re_i | ca_bus_we_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:139:50  */
  assign n1183_o = 1'b1 ? n1181_o : ca_bus_re_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:140:34  */
  assign n1184_o = cb_bus_re_i | cb_bus_we_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:140:50  */
  assign n1186_o = 1'b0 ? n1184_o : cb_bus_re_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:143:36  */
  assign n1187_o = ca_rd_req_buf | ca_wr_req_buf;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:143:54  */
  assign n1189_o = 1'b1 ? n1187_o : ca_rd_req_buf;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:144:36  */
  assign n1190_o = cb_rd_req_buf | cb_wr_req_buf;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:144:54  */
  assign n1192_o = 1'b0 ? n1190_o : cb_rd_req_buf;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:151:34  */
  assign n1194_o = arbiter[2:0];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:157:18  */
  assign n1198_o = arbiter[2:0];
  assign n1207_o = {1'b1, 3'b100};
  assign n1208_o = {1'b0, n1194_o};
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:170:9  */
  assign n1209_o = cb_req_pending ? n1207_o : n1208_o;
  assign n1210_o = {1'b1, 3'b011};
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:167:9  */
  assign n1211_o = cb_req_current ? n1210_o : n1209_o;
  assign n1212_o = {1'b0, 3'b010};
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:164:9  */
  assign n1213_o = ca_req_pending ? n1212_o : n1211_o;
  assign n1214_o = {1'b0, 3'b001};
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:161:9  */
  assign n1215_o = ca_req_current ? n1214_o : n1213_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:159:7  */
  assign n1217_o = n1198_o == 3'b000;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:178:32  */
  assign n1219_o = p_bus_err_i | p_bus_ack_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:179:37  */
  assign n1220_o = cb_req_pending | cb_req_current;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:179:11  */
  assign n1223_o = n1220_o ? 3'b100 : 3'b000;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:178:9  */
  assign n1224_o = n1219_o ? n1223_o : n1194_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:175:7  */
  assign n1226_o = n1198_o == 3'b001;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:186:7  */
  assign n1230_o = n1198_o == 3'b010;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:196:32  */
  assign n1232_o = p_bus_err_i | p_bus_ack_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:197:37  */
  assign n1233_o = ca_req_pending | ca_req_current;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:197:11  */
  assign n1236_o = n1233_o ? 3'b010 : 3'b000;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:196:9  */
  assign n1237_o = n1232_o ? n1236_o : n1194_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:193:7  */
  assign n1239_o = n1198_o == 3'b011;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:204:7  */
  assign n1243_o = n1198_o == 3'b100;
  assign n1245_o = {n1243_o, n1239_o, n1230_o, n1226_o, n1217_o};
  assign n1246_o = n1215_o[2:0];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:157:5  */
  always @*
    case (n1245_o)
      5'b10000: n1247_o = 3'b011;
      5'b01000: n1247_o = n1237_o;
      5'b00100: n1247_o = 3'b001;
      5'b00010: n1247_o = n1224_o;
      5'b00001: n1247_o = n1246_o;
      default: n1247_o = 3'b000;
    endcase
  assign n1248_o = n1215_o[3];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:157:5  */
  always @*
    case (n1245_o)
      5'b10000: n1249_o = 1'b1;
      5'b01000: n1249_o = 1'b1;
      5'b00100: n1249_o = 1'b0;
      5'b00010: n1249_o = 1'b0;
      5'b00001: n1249_o = n1248_o;
      default: n1249_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:157:5  */
  always @*
    case (n1245_o)
      5'b10000: n1250_o = cb_rd_req_buf;
      5'b01000: n1250_o = 1'b0;
      5'b00100: n1250_o = ca_rd_req_buf;
      5'b00010: n1250_o = 1'b0;
      5'b00001: n1250_o = 1'b0;
      default: n1250_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:157:5  */
  always @*
    case (n1245_o)
      5'b10000: n1251_o = cb_wr_req_buf;
      5'b01000: n1251_o = 1'b0;
      5'b00100: n1251_o = ca_wr_req_buf;
      5'b00010: n1251_o = 1'b0;
      5'b00001: n1251_o = 1'b0;
      default: n1251_o = 1'b0;
    endcase
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:221:49  */
  assign n1253_o = arbiter[6];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:221:57  */
  assign n1254_o = ~n1253_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:221:35  */
  assign n1255_o = n1254_o ? ca_bus_addr_i : cb_bus_addr_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:223:36  */
  assign n1257_o = 1'b0 ? cb_bus_wdata_i : n1259_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:223:68  */
  assign n1259_o = 1'b1 ? ca_bus_wdata_i : n1262_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:225:50  */
  assign n1260_o = arbiter[6];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:225:58  */
  assign n1261_o = ~n1260_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:224:68  */
  assign n1262_o = n1261_o ? ca_bus_wdata_i : cb_bus_wdata_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:227:34  */
  assign n1264_o = 1'b0 ? cb_bus_ben_i : n1266_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:227:66  */
  assign n1266_o = 1'b1 ? ca_bus_ben_i : n1269_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:229:48  */
  assign n1267_o = arbiter[6];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:229:56  */
  assign n1268_o = ~n1267_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:228:66  */
  assign n1269_o = n1268_o ? ca_bus_ben_i : cb_bus_ben_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:231:51  */
  assign n1270_o = arbiter[6];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:231:59  */
  assign n1271_o = ~n1270_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:231:37  */
  assign n1272_o = n1271_o ? ca_bus_cached_i : cb_bus_cached_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:232:51  */
  assign n1273_o = arbiter[6];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:232:59  */
  assign n1274_o = ~n1273_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:232:37  */
  assign n1275_o = n1274_o ? ca_bus_priv_i : cb_bus_priv_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:234:47  */
  assign n1276_o = arbiter[6];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:234:55  */
  assign n1277_o = ~n1276_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:234:33  */
  assign n1278_o = n1277_o ? ca_bus_we_i : cb_bus_we_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:235:47  */
  assign n1279_o = arbiter[6];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:235:55  */
  assign n1280_o = ~n1279_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:235:33  */
  assign n1281_o = n1280_o ? ca_bus_re_i : cb_bus_re_i;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:236:41  */
  assign n1282_o = arbiter[8];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:236:30  */
  assign n1283_o = p_bus_we | n1282_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:237:41  */
  assign n1284_o = arbiter[7];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:237:30  */
  assign n1285_o = p_bus_re | n1284_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:239:29  */
  assign n1286_o = arbiter[6];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:244:47  */
  assign n1287_o = arbiter[6];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:244:55  */
  assign n1288_o = ~n1287_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:244:33  */
  assign n1289_o = n1288_o ? p_bus_ack_i : 1'b0;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:245:47  */
  assign n1291_o = arbiter[6];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:245:33  */
  assign n1292_o = n1291_o ? p_bus_ack_i : 1'b0;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:249:47  */
  assign n1294_o = arbiter[6];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:249:55  */
  assign n1295_o = ~n1294_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:249:33  */
  assign n1296_o = n1295_o ? p_bus_err_i : 1'b0;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:250:47  */
  assign n1298_o = arbiter[6];
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:250:33  */
  assign n1299_o = n1298_o ? p_bus_err_i : 1'b0;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:127:5  */
  always @(posedge clk_i or posedge n1139_o)
    if (n1139_o)
      n1301_q <= 1'b0;
    else
      n1301_q <= n1146_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:127:5  */
  always @(posedge clk_i or posedge n1139_o)
    if (n1139_o)
      n1302_q <= 1'b0;
    else
      n1302_q <= n1153_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:127:5  */
  always @(posedge clk_i or posedge n1139_o)
    if (n1139_o)
      n1303_q <= 1'b0;
    else
      n1303_q <= n1157_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:127:5  */
  always @(posedge clk_i or posedge n1139_o)
    if (n1139_o)
      n1304_q <= 1'b0;
    else
      n1304_q <= n1164_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:127:5  */
  always @(posedge clk_i or posedge n1139_o)
    if (n1139_o)
      n1305_q <= 3'b000;
    else
      n1305_q <= n1142_o;
  /* ../neorv32/rtl/core/neorv32_busswitch.vhd:121:5  */
  assign n1306_o = {n1251_o, n1250_o, n1249_o, n1247_o, n1305_q};
endmodule

module neorv32_cpu_1_0_4_0_40_8cd82fcc1d144656bad81224642c94d0248852b6
  (input  clk_i,
   input  rstn_i,
   input  [31:0] i_bus_rdata_i,
   input  i_bus_ack_i,
   input  i_bus_err_i,
   input  [31:0] d_bus_rdata_i,
   input  d_bus_ack_i,
   input  d_bus_err_i,
   input  msw_irq_i,
   input  mext_irq_i,
   input  mtime_irq_i,
   input  [15:0] firq_i,
   input  db_halt_req_i,
   output sleep_o,
   output debug_o,
   output [31:0] i_bus_addr_o,
   output i_bus_re_o,
   output i_bus_fence_o,
   output i_bus_priv_o,
   output [31:0] d_bus_addr_o,
   output [31:0] d_bus_wdata_o,
   output [3:0] d_bus_ben_o,
   output d_bus_we_o,
   output d_bus_re_o,
   output d_bus_fence_o,
   output d_bus_priv_o);
  wire [69:0] ctrl;
  wire [31:0] imm;
  wire [31:0] rs1;
  wire [31:0] rs2;
  wire [31:0] rs3;
  wire [31:0] rs4;
  wire [31:0] alu_res;
  wire [31:0] alu_add;
  wire [1:0] alu_cmp;
  wire [31:0] mem_rdata;
  wire cp_done;
  wire alu_exc;
  wire bus_d_wait;
  wire [31:0] csr_rdata;
  wire [31:0] mar;
  wire ma_load;
  wire ma_store;
  wire be_load;
  wire be_store;
  wire [31:0] fetch_pc;
  wire [31:0] curr_pc;
  wire [31:0] next_pc;
  wire [4:0] fpu_flags;
  wire i_pmp_fault;
  wire [543:0] pmp_addr;
  wire [127:0] pmp_ctrl;
  wire [69:0] neorv32_cpu_control_inst_n942;
  wire [31:0] neorv32_cpu_control_inst_n943;
  wire neorv32_cpu_control_inst_n944;
  wire [31:0] neorv32_cpu_control_inst_n945;
  wire [31:0] neorv32_cpu_control_inst_n946;
  wire [31:0] neorv32_cpu_control_inst_n947;
  wire [31:0] neorv32_cpu_control_inst_n948;
  wire [543:0] neorv32_cpu_control_inst_n949;
  wire [127:0] neorv32_cpu_control_inst_n950;
  wire neorv32_cpu_control_inst_ctrl_o_rf_wb_en;
  wire [4:0] neorv32_cpu_control_inst_ctrl_o_rf_rs1;
  wire [4:0] neorv32_cpu_control_inst_ctrl_o_rf_rs2;
  wire [4:0] neorv32_cpu_control_inst_ctrl_o_rf_rs3;
  wire [4:0] neorv32_cpu_control_inst_ctrl_o_rf_rd;
  wire [1:0] neorv32_cpu_control_inst_ctrl_o_rf_mux;
  wire neorv32_cpu_control_inst_ctrl_o_rf_zero_we;
  wire [2:0] neorv32_cpu_control_inst_ctrl_o_alu_op;
  wire neorv32_cpu_control_inst_ctrl_o_alu_opa_mux;
  wire neorv32_cpu_control_inst_ctrl_o_alu_opb_mux;
  wire neorv32_cpu_control_inst_ctrl_o_alu_unsigned;
  wire [2:0] neorv32_cpu_control_inst_ctrl_o_alu_frm;
  wire [5:0] neorv32_cpu_control_inst_ctrl_o_alu_cp_trig;
  wire neorv32_cpu_control_inst_ctrl_o_bus_req;
  wire neorv32_cpu_control_inst_ctrl_o_bus_mo_we;
  wire neorv32_cpu_control_inst_ctrl_o_bus_fence;
  wire neorv32_cpu_control_inst_ctrl_o_bus_fencei;
  wire neorv32_cpu_control_inst_ctrl_o_bus_priv;
  wire [2:0] neorv32_cpu_control_inst_ctrl_o_ir_funct3;
  wire [11:0] neorv32_cpu_control_inst_ctrl_o_ir_funct12;
  wire [6:0] neorv32_cpu_control_inst_ctrl_o_ir_opcode;
  wire neorv32_cpu_control_inst_ctrl_o_cpu_priv;
  wire neorv32_cpu_control_inst_ctrl_o_cpu_sleep;
  wire neorv32_cpu_control_inst_ctrl_o_cpu_trap;
  wire neorv32_cpu_control_inst_ctrl_o_cpu_debug;
  wire [31:0] neorv32_cpu_control_inst_i_bus_addr_o;
  wire neorv32_cpu_control_inst_i_bus_re_o;
  wire [31:0] neorv32_cpu_control_inst_imm_o;
  wire [31:0] neorv32_cpu_control_inst_curr_pc_o;
  wire [31:0] neorv32_cpu_control_inst_next_pc_o;
  wire [31:0] neorv32_cpu_control_inst_csr_rdata_o;
  wire [543:0] neorv32_cpu_control_inst_pmp_addr_o;
  wire [127:0] neorv32_cpu_control_inst_pmp_ctrl_o;
  wire [69:0] n951_o;
  wire n970_o;
  wire n971_o;
  wire n972_o;
  wire n973_o;
  wire [31:0] neorv32_cpu_regfile_inst_n974;
  wire [31:0] neorv32_cpu_regfile_inst_n975;
  wire [31:0] neorv32_cpu_regfile_inst_n976;
  wire [31:0] neorv32_cpu_regfile_inst_n977;
  wire [31:0] neorv32_cpu_regfile_inst_rs1_o;
  wire [31:0] neorv32_cpu_regfile_inst_rs2_o;
  wire [31:0] neorv32_cpu_regfile_inst_rs3_o;
  wire [31:0] neorv32_cpu_regfile_inst_rs4_o;
  wire n978_o;
  wire [4:0] n979_o;
  wire [4:0] n980_o;
  wire [4:0] n981_o;
  wire [4:0] n982_o;
  wire [1:0] n983_o;
  wire n984_o;
  wire [2:0] n985_o;
  wire n986_o;
  wire n987_o;
  wire n988_o;
  wire [2:0] n989_o;
  wire [5:0] n990_o;
  wire n991_o;
  wire n992_o;
  wire n993_o;
  wire n994_o;
  wire n995_o;
  wire [2:0] n996_o;
  wire [11:0] n997_o;
  wire [6:0] n998_o;
  wire n999_o;
  wire n1000_o;
  wire n1001_o;
  wire n1002_o;
  wire [1:0] neorv32_cpu_alu_inst_n1011;
  wire [31:0] neorv32_cpu_alu_inst_n1012;
  wire [31:0] neorv32_cpu_alu_inst_n1013;
  wire [4:0] neorv32_cpu_alu_inst_n1014;
  wire neorv32_cpu_alu_inst_n1015;
  wire neorv32_cpu_alu_inst_n1016;
  wire [1:0] neorv32_cpu_alu_inst_cmp_o;
  wire [31:0] neorv32_cpu_alu_inst_res_o;
  wire [31:0] neorv32_cpu_alu_inst_add_o;
  wire [4:0] neorv32_cpu_alu_inst_fpu_flags_o;
  wire neorv32_cpu_alu_inst_exc_o;
  wire neorv32_cpu_alu_inst_cp_done_o;
  wire n1017_o;
  wire [4:0] n1018_o;
  wire [4:0] n1019_o;
  wire [4:0] n1020_o;
  wire [4:0] n1021_o;
  wire [1:0] n1022_o;
  wire n1023_o;
  wire [2:0] n1024_o;
  wire n1025_o;
  wire n1026_o;
  wire n1027_o;
  wire [2:0] n1028_o;
  wire [5:0] n1029_o;
  wire n1030_o;
  wire n1031_o;
  wire n1032_o;
  wire n1033_o;
  wire n1034_o;
  wire [2:0] n1035_o;
  wire [11:0] n1036_o;
  wire [6:0] n1037_o;
  wire n1038_o;
  wire n1039_o;
  wire n1040_o;
  wire n1041_o;
  wire neorv32_cpu_bus_inst_n1054;
  wire [31:0] neorv32_cpu_bus_inst_n1055;
  wire [31:0] neorv32_cpu_bus_inst_n1056;
  wire neorv32_cpu_bus_inst_n1057;
  wire neorv32_cpu_bus_inst_n1058;
  wire neorv32_cpu_bus_inst_n1059;
  wire neorv32_cpu_bus_inst_n1060;
  wire neorv32_cpu_bus_inst_n1061;
  wire [31:0] neorv32_cpu_bus_inst_n1062;
  wire [31:0] neorv32_cpu_bus_inst_n1063;
  wire [3:0] neorv32_cpu_bus_inst_n1064;
  wire neorv32_cpu_bus_inst_n1065;
  wire neorv32_cpu_bus_inst_n1066;
  wire neorv32_cpu_bus_inst_n1067;
  wire neorv32_cpu_bus_inst_n1068;
  wire neorv32_cpu_bus_inst_i_pmp_fault_o;
  wire [31:0] neorv32_cpu_bus_inst_rdata_o;
  wire [31:0] neorv32_cpu_bus_inst_mar_o;
  wire neorv32_cpu_bus_inst_d_wait_o;
  wire neorv32_cpu_bus_inst_ma_load_o;
  wire neorv32_cpu_bus_inst_ma_store_o;
  wire neorv32_cpu_bus_inst_be_load_o;
  wire neorv32_cpu_bus_inst_be_store_o;
  wire [31:0] neorv32_cpu_bus_inst_d_bus_addr_o;
  wire [31:0] neorv32_cpu_bus_inst_d_bus_wdata_o;
  wire [3:0] neorv32_cpu_bus_inst_d_bus_ben_o;
  wire neorv32_cpu_bus_inst_d_bus_we_o;
  wire neorv32_cpu_bus_inst_d_bus_re_o;
  wire neorv32_cpu_bus_inst_d_bus_fence_o;
  wire neorv32_cpu_bus_inst_d_bus_priv_o;
  wire n1069_o;
  wire [4:0] n1070_o;
  wire [4:0] n1071_o;
  wire [4:0] n1072_o;
  wire [4:0] n1073_o;
  wire [1:0] n1074_o;
  wire n1075_o;
  wire [2:0] n1076_o;
  wire n1077_o;
  wire n1078_o;
  wire n1079_o;
  wire [2:0] n1080_o;
  wire [5:0] n1081_o;
  wire n1082_o;
  wire n1083_o;
  wire n1084_o;
  wire n1085_o;
  wire n1086_o;
  wire [2:0] n1087_o;
  wire [11:0] n1088_o;
  wire [6:0] n1089_o;
  wire n1090_o;
  wire n1091_o;
  wire n1092_o;
  wire n1093_o;
  assign sleep_o = n970_o;
  assign debug_o = n971_o;
  assign i_bus_addr_o = fetch_pc;
  assign i_bus_re_o = neorv32_cpu_control_inst_n944;
  assign i_bus_fence_o = n972_o;
  assign i_bus_priv_o = n973_o;
  assign d_bus_addr_o = neorv32_cpu_bus_inst_n1062;
  assign d_bus_wdata_o = neorv32_cpu_bus_inst_n1063;
  assign d_bus_ben_o = neorv32_cpu_bus_inst_n1064;
  assign d_bus_we_o = neorv32_cpu_bus_inst_n1065;
  assign d_bus_re_o = neorv32_cpu_bus_inst_n1066;
  assign d_bus_fence_o = neorv32_cpu_bus_inst_n1067;
  assign d_bus_priv_o = neorv32_cpu_bus_inst_n1068;
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:128:10  */
  assign ctrl = neorv32_cpu_control_inst_n942; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:129:10  */
  assign imm = neorv32_cpu_control_inst_n945; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:130:10  */
  assign rs1 = neorv32_cpu_regfile_inst_n974; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:131:10  */
  assign rs2 = neorv32_cpu_regfile_inst_n975; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:132:10  */
  assign rs3 = neorv32_cpu_regfile_inst_n976; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:133:10  */
  assign rs4 = neorv32_cpu_regfile_inst_n977; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:134:10  */
  assign alu_res = neorv32_cpu_alu_inst_n1012; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:135:10  */
  assign alu_add = neorv32_cpu_alu_inst_n1013; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:136:10  */
  assign alu_cmp = neorv32_cpu_alu_inst_n1011; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:137:10  */
  assign mem_rdata = neorv32_cpu_bus_inst_n1055; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:138:10  */
  assign cp_done = neorv32_cpu_alu_inst_n1016; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:139:10  */
  assign alu_exc = neorv32_cpu_alu_inst_n1015; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:140:10  */
  assign bus_d_wait = neorv32_cpu_bus_inst_n1057; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:141:10  */
  assign csr_rdata = neorv32_cpu_control_inst_n948; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:142:10  */
  assign mar = neorv32_cpu_bus_inst_n1056; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:143:10  */
  assign ma_load = neorv32_cpu_bus_inst_n1058; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:144:10  */
  assign ma_store = neorv32_cpu_bus_inst_n1059; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:145:10  */
  assign be_load = neorv32_cpu_bus_inst_n1060; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:146:10  */
  assign be_store = neorv32_cpu_bus_inst_n1061; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:147:10  */
  assign fetch_pc = neorv32_cpu_control_inst_n943; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:148:10  */
  assign curr_pc = neorv32_cpu_control_inst_n946; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:149:10  */
  assign next_pc = neorv32_cpu_control_inst_n947; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:150:10  */
  assign fpu_flags = neorv32_cpu_alu_inst_n1014; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:151:10  */
  assign i_pmp_fault = neorv32_cpu_bus_inst_n1054; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:154:10  */
  assign pmp_addr = neorv32_cpu_control_inst_n949; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:155:10  */
  assign pmp_ctrl = neorv32_cpu_control_inst_n950; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:280:22  */
  assign neorv32_cpu_control_inst_n942 = n951_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:282:22  */
  assign neorv32_cpu_control_inst_n943 = neorv32_cpu_control_inst_i_bus_addr_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:284:22  */
  assign neorv32_cpu_control_inst_n944 = neorv32_cpu_control_inst_i_bus_re_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:297:22  */
  assign neorv32_cpu_control_inst_n945 = neorv32_cpu_control_inst_imm_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:298:22  */
  assign neorv32_cpu_control_inst_n946 = neorv32_cpu_control_inst_curr_pc_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:299:22  */
  assign neorv32_cpu_control_inst_n947 = neorv32_cpu_control_inst_next_pc_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:300:22  */
  assign neorv32_cpu_control_inst_n948 = neorv32_cpu_control_inst_csr_rdata_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:312:22  */
  assign neorv32_cpu_control_inst_n949 = neorv32_cpu_control_inst_pmp_addr_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:313:22  */
  assign neorv32_cpu_control_inst_n950 = neorv32_cpu_control_inst_pmp_ctrl_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:241:3  */
  neorv32_cpu_control_32_2_0_4_0_40_8cd82fcc1d144656bad81224642c94d0248852b6 neorv32_cpu_control_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .i_bus_rdata_i(i_bus_rdata_i),
    .i_bus_ack_i(i_bus_ack_i),
    .i_bus_err_i(i_bus_err_i),
    .i_pmp_fault_i(i_pmp_fault),
    .alu_cp_done_i(cp_done),
    .alu_exc_i(alu_exc),
    .bus_d_wait_i(bus_d_wait),
    .cmp_i(alu_cmp),
    .alu_add_i(alu_add),
    .rs1_i(rs1),
    .fpu_flags_i(fpu_flags),
    .db_halt_req_i(db_halt_req_i),
    .msw_irq_i(msw_irq_i),
    .mext_irq_i(mext_irq_i),
    .mtime_irq_i(mtime_irq_i),
    .firq_i(firq_i),
    .mar_i(mar),
    .ma_load_i(ma_load),
    .ma_store_i(ma_store),
    .be_load_i(be_load),
    .be_store_i(be_store),
    .ctrl_o_rf_wb_en(neorv32_cpu_control_inst_ctrl_o_rf_wb_en),
    .ctrl_o_rf_rs1(neorv32_cpu_control_inst_ctrl_o_rf_rs1),
    .ctrl_o_rf_rs2(neorv32_cpu_control_inst_ctrl_o_rf_rs2),
    .ctrl_o_rf_rs3(neorv32_cpu_control_inst_ctrl_o_rf_rs3),
    .ctrl_o_rf_rd(neorv32_cpu_control_inst_ctrl_o_rf_rd),
    .ctrl_o_rf_mux(neorv32_cpu_control_inst_ctrl_o_rf_mux),
    .ctrl_o_rf_zero_we(neorv32_cpu_control_inst_ctrl_o_rf_zero_we),
    .ctrl_o_alu_op(neorv32_cpu_control_inst_ctrl_o_alu_op),
    .ctrl_o_alu_opa_mux(neorv32_cpu_control_inst_ctrl_o_alu_opa_mux),
    .ctrl_o_alu_opb_mux(neorv32_cpu_control_inst_ctrl_o_alu_opb_mux),
    .ctrl_o_alu_unsigned(neorv32_cpu_control_inst_ctrl_o_alu_unsigned),
    .ctrl_o_alu_frm(neorv32_cpu_control_inst_ctrl_o_alu_frm),
    .ctrl_o_alu_cp_trig(neorv32_cpu_control_inst_ctrl_o_alu_cp_trig),
    .ctrl_o_bus_req(neorv32_cpu_control_inst_ctrl_o_bus_req),
    .ctrl_o_bus_mo_we(neorv32_cpu_control_inst_ctrl_o_bus_mo_we),
    .ctrl_o_bus_fence(neorv32_cpu_control_inst_ctrl_o_bus_fence),
    .ctrl_o_bus_fencei(neorv32_cpu_control_inst_ctrl_o_bus_fencei),
    .ctrl_o_bus_priv(neorv32_cpu_control_inst_ctrl_o_bus_priv),
    .ctrl_o_ir_funct3(neorv32_cpu_control_inst_ctrl_o_ir_funct3),
    .ctrl_o_ir_funct12(neorv32_cpu_control_inst_ctrl_o_ir_funct12),
    .ctrl_o_ir_opcode(neorv32_cpu_control_inst_ctrl_o_ir_opcode),
    .ctrl_o_cpu_priv(neorv32_cpu_control_inst_ctrl_o_cpu_priv),
    .ctrl_o_cpu_sleep(neorv32_cpu_control_inst_ctrl_o_cpu_sleep),
    .ctrl_o_cpu_trap(neorv32_cpu_control_inst_ctrl_o_cpu_trap),
    .ctrl_o_cpu_debug(neorv32_cpu_control_inst_ctrl_o_cpu_debug),
    .i_bus_addr_o(neorv32_cpu_control_inst_i_bus_addr_o),
    .i_bus_re_o(neorv32_cpu_control_inst_i_bus_re_o),
    .imm_o(neorv32_cpu_control_inst_imm_o),
    .curr_pc_o(neorv32_cpu_control_inst_curr_pc_o),
    .next_pc_o(neorv32_cpu_control_inst_next_pc_o),
    .csr_rdata_o(neorv32_cpu_control_inst_csr_rdata_o),
    .pmp_addr_o(neorv32_cpu_control_inst_pmp_addr_o),
    .pmp_ctrl_o(neorv32_cpu_control_inst_pmp_ctrl_o));
  /* ../neorv32/rtl/core/neorv32_top.vhd:890:17  */
  assign n951_o = {neorv32_cpu_control_inst_ctrl_o_cpu_debug, neorv32_cpu_control_inst_ctrl_o_cpu_trap, neorv32_cpu_control_inst_ctrl_o_cpu_sleep, neorv32_cpu_control_inst_ctrl_o_cpu_priv, neorv32_cpu_control_inst_ctrl_o_ir_opcode, neorv32_cpu_control_inst_ctrl_o_ir_funct12, neorv32_cpu_control_inst_ctrl_o_ir_funct3, neorv32_cpu_control_inst_ctrl_o_bus_priv, neorv32_cpu_control_inst_ctrl_o_bus_fencei, neorv32_cpu_control_inst_ctrl_o_bus_fence, neorv32_cpu_control_inst_ctrl_o_bus_mo_we, neorv32_cpu_control_inst_ctrl_o_bus_req, neorv32_cpu_control_inst_ctrl_o_alu_cp_trig, neorv32_cpu_control_inst_ctrl_o_alu_frm, neorv32_cpu_control_inst_ctrl_o_alu_unsigned, neorv32_cpu_control_inst_ctrl_o_alu_opb_mux, neorv32_cpu_control_inst_ctrl_o_alu_opa_mux, neorv32_cpu_control_inst_ctrl_o_alu_op, neorv32_cpu_control_inst_ctrl_o_rf_zero_we, neorv32_cpu_control_inst_ctrl_o_rf_mux, neorv32_cpu_control_inst_ctrl_o_rf_rd, neorv32_cpu_control_inst_ctrl_o_rf_rs3, neorv32_cpu_control_inst_ctrl_o_rf_rs2, neorv32_cpu_control_inst_ctrl_o_rf_rs1, neorv32_cpu_control_inst_ctrl_o_rf_wb_en};
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:323:19  */
  assign n970_o = ctrl[67];
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:324:19  */
  assign n971_o = ctrl[69];
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:328:25  */
  assign n972_o = ctrl[42];
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:329:25  */
  assign n973_o = ctrl[66];
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:351:15  */
  assign neorv32_cpu_regfile_inst_n974 = neorv32_cpu_regfile_inst_rs1_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:352:15  */
  assign neorv32_cpu_regfile_inst_n975 = neorv32_cpu_regfile_inst_rs2_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:353:15  */
  assign neorv32_cpu_regfile_inst_n976 = neorv32_cpu_regfile_inst_rs3_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:354:15  */
  assign neorv32_cpu_regfile_inst_n977 = neorv32_cpu_regfile_inst_rs4_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:334:3  */
  neorv32_cpu_regfile_32_29e2dcfbb16f63bb0254df7585a15bb6fb5e927d neorv32_cpu_regfile_inst (
    .clk_i(clk_i),
    .ctrl_i_rf_wb_en(n978_o),
    .ctrl_i_rf_rs1(n979_o),
    .ctrl_i_rf_rs2(n980_o),
    .ctrl_i_rf_rs3(n981_o),
    .ctrl_i_rf_rd(n982_o),
    .ctrl_i_rf_mux(n983_o),
    .ctrl_i_rf_zero_we(n984_o),
    .ctrl_i_alu_op(n985_o),
    .ctrl_i_alu_opa_mux(n986_o),
    .ctrl_i_alu_opb_mux(n987_o),
    .ctrl_i_alu_unsigned(n988_o),
    .ctrl_i_alu_frm(n989_o),
    .ctrl_i_alu_cp_trig(n990_o),
    .ctrl_i_bus_req(n991_o),
    .ctrl_i_bus_mo_we(n992_o),
    .ctrl_i_bus_fence(n993_o),
    .ctrl_i_bus_fencei(n994_o),
    .ctrl_i_bus_priv(n995_o),
    .ctrl_i_ir_funct3(n996_o),
    .ctrl_i_ir_funct12(n997_o),
    .ctrl_i_ir_opcode(n998_o),
    .ctrl_i_cpu_priv(n999_o),
    .ctrl_i_cpu_sleep(n1000_o),
    .ctrl_i_cpu_trap(n1001_o),
    .ctrl_i_cpu_debug(n1002_o),
    .alu_i(alu_res),
    .mem_i(mem_rdata),
    .csr_i(csr_rdata),
    .pc2_i(next_pc),
    .rs1_o(neorv32_cpu_regfile_inst_rs1_o),
    .rs2_o(neorv32_cpu_regfile_inst_rs2_o),
    .rs3_o(neorv32_cpu_regfile_inst_rs3_o),
    .rs4_o(neorv32_cpu_regfile_inst_rs4_o));
  /* ../neorv32/rtl/core/neorv32_top.vhd:748:24  */
  assign n978_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:747:24  */
  assign n979_o = ctrl[5:1];
  /* ../neorv32/rtl/core/neorv32_top.vhd:745:24  */
  assign n980_o = ctrl[10:6];
  /* ../neorv32/rtl/core/neorv32_top.vhd:744:24  */
  assign n981_o = ctrl[15:11];
  /* ../neorv32/rtl/core/neorv32_top.vhd:739:24  */
  assign n982_o = ctrl[20:16];
  /* ../neorv32/rtl/core/neorv32_top.vhd:734:24  */
  assign n983_o = ctrl[22:21];
  /* ../neorv32/rtl/core/neorv32_top.vhd:733:24  */
  assign n984_o = ctrl[23];
  /* ../neorv32/rtl/core/neorv32_top.vhd:728:24  */
  assign n985_o = ctrl[26:24];
  /* ../neorv32/rtl/core/neorv32_top.vhd:715:3  */
  assign n986_o = ctrl[27];
  /* ../neorv32/rtl/core/neorv32_top.vhd:715:3  */
  assign n987_o = ctrl[28];
  /* ../neorv32/rtl/core/neorv32_top.vhd:715:3  */
  assign n988_o = ctrl[29];
  /* ../neorv32/rtl/core/neorv32_top.vhd:715:3  */
  assign n989_o = ctrl[32:30];
  /* ../neorv32/rtl/core/neorv32_top.vhd:715:3  */
  assign n990_o = ctrl[38:33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:715:3  */
  assign n991_o = ctrl[39];
  /* ../neorv32/rtl/core/neorv32_top.vhd:715:3  */
  assign n992_o = ctrl[40];
  /* ../neorv32/rtl/core/neorv32_top.vhd:715:3  */
  assign n993_o = ctrl[41];
  /* ../neorv32/rtl/core/neorv32_top.vhd:715:3  */
  assign n994_o = ctrl[42];
  /* ../neorv32/rtl/core/neorv32_top.vhd:715:3  */
  assign n995_o = ctrl[43];
  /* ../neorv32/rtl/core/neorv32_top.vhd:715:3  */
  assign n996_o = ctrl[46:44];
  /* ../neorv32/rtl/core/neorv32_top.vhd:715:3  */
  assign n997_o = ctrl[58:47];
  /* ../neorv32/rtl/core/neorv32_top.vhd:715:3  */
  assign n998_o = ctrl[65:59];
  /* ../neorv32/rtl/core/neorv32_top.vhd:715:3  */
  assign n999_o = ctrl[66];
  /* ../neorv32/rtl/core/neorv32_top.vhd:572:22  */
  assign n1000_o = ctrl[67];
  /* ../neorv32/rtl/core/neorv32_top.vhd:571:22  */
  assign n1001_o = ctrl[68];
  /* ../neorv32/rtl/core/neorv32_top.vhd:568:22  */
  assign n1002_o = ctrl[69];
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:387:20  */
  assign neorv32_cpu_alu_inst_n1011 = neorv32_cpu_alu_inst_cmp_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:388:20  */
  assign neorv32_cpu_alu_inst_n1012 = neorv32_cpu_alu_inst_res_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:389:20  */
  assign neorv32_cpu_alu_inst_n1013 = neorv32_cpu_alu_inst_add_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:390:20  */
  assign neorv32_cpu_alu_inst_n1014 = neorv32_cpu_alu_inst_fpu_flags_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:392:20  */
  assign neorv32_cpu_alu_inst_n1015 = neorv32_cpu_alu_inst_exc_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:393:20  */
  assign neorv32_cpu_alu_inst_n1016 = neorv32_cpu_alu_inst_cp_done_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:360:3  */
  neorv32_cpu_alu_32_5e99b7dbd159708117122aa5c1c1bfccec006ed0 neorv32_cpu_alu_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .ctrl_i_rf_wb_en(n1017_o),
    .ctrl_i_rf_rs1(n1018_o),
    .ctrl_i_rf_rs2(n1019_o),
    .ctrl_i_rf_rs3(n1020_o),
    .ctrl_i_rf_rd(n1021_o),
    .ctrl_i_rf_mux(n1022_o),
    .ctrl_i_rf_zero_we(n1023_o),
    .ctrl_i_alu_op(n1024_o),
    .ctrl_i_alu_opa_mux(n1025_o),
    .ctrl_i_alu_opb_mux(n1026_o),
    .ctrl_i_alu_unsigned(n1027_o),
    .ctrl_i_alu_frm(n1028_o),
    .ctrl_i_alu_cp_trig(n1029_o),
    .ctrl_i_bus_req(n1030_o),
    .ctrl_i_bus_mo_we(n1031_o),
    .ctrl_i_bus_fence(n1032_o),
    .ctrl_i_bus_fencei(n1033_o),
    .ctrl_i_bus_priv(n1034_o),
    .ctrl_i_ir_funct3(n1035_o),
    .ctrl_i_ir_funct12(n1036_o),
    .ctrl_i_ir_opcode(n1037_o),
    .ctrl_i_cpu_priv(n1038_o),
    .ctrl_i_cpu_sleep(n1039_o),
    .ctrl_i_cpu_trap(n1040_o),
    .ctrl_i_cpu_debug(n1041_o),
    .rs1_i(rs1),
    .rs2_i(rs2),
    .rs3_i(rs3),
    .rs4_i(rs4),
    .pc_i(curr_pc),
    .imm_i(imm),
    .cmp_o(neorv32_cpu_alu_inst_cmp_o),
    .res_o(neorv32_cpu_alu_inst_res_o),
    .add_o(neorv32_cpu_alu_inst_add_o),
    .fpu_flags_o(neorv32_cpu_alu_inst_fpu_flags_o),
    .exc_o(neorv32_cpu_alu_inst_exc_o),
    .cp_done_o(neorv32_cpu_alu_inst_cp_done_o));
  /* ../neorv32/rtl/core/neorv32_top.vhd:514:3  */
  assign n1017_o = ctrl[0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:514:3  */
  assign n1018_o = ctrl[5:1];
  /* ../neorv32/rtl/core/neorv32_top.vhd:514:3  */
  assign n1019_o = ctrl[10:6];
  /* ../neorv32/rtl/core/neorv32_top.vhd:514:3  */
  assign n1020_o = ctrl[15:11];
  /* ../neorv32/rtl/core/neorv32_top.vhd:226:5  */
  assign n1021_o = ctrl[20:16];
  /* ../neorv32/rtl/core/neorv32_top.vhd:223:5  */
  assign n1022_o = ctrl[22:21];
  /* ../neorv32/rtl/core/neorv32_top.vhd:219:5  */
  assign n1023_o = ctrl[23];
  /* ../neorv32/rtl/core/neorv32_top.vhd:216:5  */
  assign n1024_o = ctrl[26:24];
  /* ../neorv32/rtl/core/neorv32_top.vhd:212:5  */
  assign n1025_o = ctrl[27];
  /* ../neorv32/rtl/core/neorv32_top.vhd:210:5  */
  assign n1026_o = ctrl[28];
  /* ../neorv32/rtl/core/neorv32_top.vhd:204:5  */
  assign n1027_o = ctrl[29];
  /* ../neorv32/rtl/core/neorv32_top.vhd:200:5  */
  assign n1028_o = ctrl[32:30];
  /* ../neorv32/rtl/core/neorv32_top.vhd:198:5  */
  assign n1029_o = ctrl[38:33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:197:5  */
  assign n1030_o = ctrl[39];
  /* ../neorv32/rtl/core/neorv32_top.vhd:193:5  */
  assign n1031_o = ctrl[40];
  /* ../neorv32/rtl/core/neorv32_top.vhd:191:5  */
  assign n1032_o = ctrl[41];
  /* ../neorv32/rtl/core/neorv32_top.vhd:187:5  */
  assign n1033_o = ctrl[42];
  /* ../neorv32/rtl/core/neorv32_top.vhd:185:5  */
  assign n1034_o = ctrl[43];
  /* ../neorv32/rtl/core/neorv32_top.vhd:181:5  */
  assign n1035_o = ctrl[46:44];
  /* ../neorv32/rtl/core/neorv32_top.vhd:178:5  */
  assign n1036_o = ctrl[58:47];
  /* ../neorv32/rtl/core/neorv32_top.vhd:176:5  */
  assign n1037_o = ctrl[65:59];
  /* ../neorv32/rtl/core/neorv32_top.vhd:175:5  */
  assign n1038_o = ctrl[66];
  /* ../neorv32/rtl/core/neorv32_top.vhd:172:5  */
  assign n1039_o = ctrl[67];
  /* ../neorv32/rtl/core/neorv32_top.vhd:171:5  */
  assign n1040_o = ctrl[68];
  /* ../neorv32/rtl/core/neorv32_top.vhd:166:5  */
  assign n1041_o = ctrl[69];
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:412:22  */
  assign neorv32_cpu_bus_inst_n1054 = neorv32_cpu_bus_inst_i_pmp_fault_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:416:22  */
  assign neorv32_cpu_bus_inst_n1055 = neorv32_cpu_bus_inst_rdata_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:417:22  */
  assign neorv32_cpu_bus_inst_n1056 = neorv32_cpu_bus_inst_mar_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:418:22  */
  assign neorv32_cpu_bus_inst_n1057 = neorv32_cpu_bus_inst_d_wait_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:419:22  */
  assign neorv32_cpu_bus_inst_n1058 = neorv32_cpu_bus_inst_ma_load_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:420:22  */
  assign neorv32_cpu_bus_inst_n1059 = neorv32_cpu_bus_inst_ma_store_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:421:22  */
  assign neorv32_cpu_bus_inst_n1060 = neorv32_cpu_bus_inst_be_load_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:422:22  */
  assign neorv32_cpu_bus_inst_n1061 = neorv32_cpu_bus_inst_be_store_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:427:22  */
  assign neorv32_cpu_bus_inst_n1062 = neorv32_cpu_bus_inst_d_bus_addr_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:429:22  */
  assign neorv32_cpu_bus_inst_n1063 = neorv32_cpu_bus_inst_d_bus_wdata_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:430:22  */
  assign neorv32_cpu_bus_inst_n1064 = neorv32_cpu_bus_inst_d_bus_ben_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:431:22  */
  assign neorv32_cpu_bus_inst_n1065 = neorv32_cpu_bus_inst_d_bus_we_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:432:22  */
  assign neorv32_cpu_bus_inst_n1066 = neorv32_cpu_bus_inst_d_bus_re_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:435:22  */
  assign neorv32_cpu_bus_inst_n1067 = neorv32_cpu_bus_inst_d_bus_fence_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:436:22  */
  assign neorv32_cpu_bus_inst_n1068 = neorv32_cpu_bus_inst_d_bus_priv_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_cpu.vhd:399:3  */
  neorv32_cpu_bus_32_0_4 neorv32_cpu_bus_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .ctrl_i_rf_wb_en(n1069_o),
    .ctrl_i_rf_rs1(n1070_o),
    .ctrl_i_rf_rs2(n1071_o),
    .ctrl_i_rf_rs3(n1072_o),
    .ctrl_i_rf_rd(n1073_o),
    .ctrl_i_rf_mux(n1074_o),
    .ctrl_i_rf_zero_we(n1075_o),
    .ctrl_i_alu_op(n1076_o),
    .ctrl_i_alu_opa_mux(n1077_o),
    .ctrl_i_alu_opb_mux(n1078_o),
    .ctrl_i_alu_unsigned(n1079_o),
    .ctrl_i_alu_frm(n1080_o),
    .ctrl_i_alu_cp_trig(n1081_o),
    .ctrl_i_bus_req(n1082_o),
    .ctrl_i_bus_mo_we(n1083_o),
    .ctrl_i_bus_fence(n1084_o),
    .ctrl_i_bus_fencei(n1085_o),
    .ctrl_i_bus_priv(n1086_o),
    .ctrl_i_ir_funct3(n1087_o),
    .ctrl_i_ir_funct12(n1088_o),
    .ctrl_i_ir_opcode(n1089_o),
    .ctrl_i_cpu_priv(n1090_o),
    .ctrl_i_cpu_sleep(n1091_o),
    .ctrl_i_cpu_trap(n1092_o),
    .ctrl_i_cpu_debug(n1093_o),
    .fetch_pc_i(fetch_pc),
    .addr_i(alu_add),
    .wdata_i(rs2),
    .pmp_addr_i(pmp_addr),
    .pmp_ctrl_i(pmp_ctrl),
    .d_bus_rdata_i(d_bus_rdata_i),
    .d_bus_ack_i(d_bus_ack_i),
    .d_bus_err_i(d_bus_err_i),
    .i_pmp_fault_o(neorv32_cpu_bus_inst_i_pmp_fault_o),
    .rdata_o(neorv32_cpu_bus_inst_rdata_o),
    .mar_o(neorv32_cpu_bus_inst_mar_o),
    .d_wait_o(neorv32_cpu_bus_inst_d_wait_o),
    .ma_load_o(neorv32_cpu_bus_inst_ma_load_o),
    .ma_store_o(neorv32_cpu_bus_inst_ma_store_o),
    .be_load_o(neorv32_cpu_bus_inst_be_load_o),
    .be_store_o(neorv32_cpu_bus_inst_be_store_o),
    .d_bus_addr_o(neorv32_cpu_bus_inst_d_bus_addr_o),
    .d_bus_wdata_o(neorv32_cpu_bus_inst_d_bus_wdata_o),
    .d_bus_ben_o(neorv32_cpu_bus_inst_d_bus_ben_o),
    .d_bus_we_o(neorv32_cpu_bus_inst_d_bus_we_o),
    .d_bus_re_o(neorv32_cpu_bus_inst_d_bus_re_o),
    .d_bus_fence_o(neorv32_cpu_bus_inst_d_bus_fence_o),
    .d_bus_priv_o(neorv32_cpu_bus_inst_d_bus_priv_o));
  assign n1069_o = ctrl[0];
  assign n1070_o = ctrl[5:1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2438:14  */
  assign n1071_o = ctrl[10:6];
  assign n1072_o = ctrl[15:11];
  /* ../neorv32/rtl/core/neorv32_package.vhd:105:12  */
  assign n1073_o = ctrl[20:16];
  /* ../neorv32/rtl/core/neorv32_package.vhd:105:12  */
  assign n1074_o = ctrl[22:21];
  assign n1075_o = ctrl[23];
  /* ../neorv32/rtl/core/neorv32_package.vhd:105:12  */
  assign n1076_o = ctrl[26:24];
  /* ../neorv32/rtl/core/neorv32_top.vhd:467:3  */
  assign n1077_o = ctrl[27];
  assign n1078_o = ctrl[28];
  assign n1079_o = ctrl[29];
  assign n1080_o = ctrl[32:30];
  assign n1081_o = ctrl[38:33];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2450:14  */
  assign n1082_o = ctrl[39];
  assign n1083_o = ctrl[40];
  /* ../neorv32/rtl/core/neorv32_package.vhd:106:12  */
  assign n1084_o = ctrl[41];
  /* ../neorv32/rtl/core/neorv32_package.vhd:106:12  */
  assign n1085_o = ctrl[42];
  assign n1086_o = ctrl[43];
  /* ../neorv32/rtl/core/neorv32_package.vhd:106:12  */
  assign n1087_o = ctrl[46:44];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2454:22  */
  assign n1088_o = ctrl[58:47];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2454:27  */
  assign n1089_o = ctrl[65:59];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2454:22  */
  assign n1090_o = ctrl[66];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2454:27  */
  assign n1091_o = ctrl[67];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2454:22  */
  assign n1092_o = ctrl[68];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2454:27  */
  assign n1093_o = ctrl[69];
endmodule

module neorv32_top_5000000_1_0_4_0_40_1024_2048_4_64_1_4_64_255_0_0_256_256_1_1_1_0_0_1_32_32_1_69ad7886168de6916fb842204ba7129434750df3
  (input  clk_i,
   input  rstn_i,
   input  jtag_trst_i,
   input  jtag_tck_i,
   input  jtag_tdi_i,
   input  jtag_tms_i,
   input  [31:0] wb_dat_i,
   input  wb_ack_i,
   input  wb_err_i,
   input  xip_dat_i,
   input  [63:0] gpio_i,
   input  uart0_rxd_i,
   input  uart0_cts_i,
   input  uart1_rxd_i,
   input  uart1_cts_i,
   input  spi_dat_i,
   input  sdi_clk_i,
   input  sdi_dat_i,
   input  sdi_csn_i,
   input  twi_sda_i,
   input  twi_scl_i,
   input  onewire_i,
   input  [31:0] cfs_in_i,
   input  [31:0] xirq_i,
   input  mtime_irq_i,
   input  msw_irq_i,
   input  mext_irq_i,
   output jtag_tdo_o,
   output [2:0] wb_tag_o,
   output [31:0] wb_adr_o,
   output [31:0] wb_dat_o,
   output wb_we_o,
   output [3:0] wb_sel_o,
   output wb_stb_o,
   output wb_cyc_o,
   output fence_o,
   output fencei_o,
   output xip_csn_o,
   output xip_clk_o,
   output xip_dat_o,
   output [63:0] gpio_o,
   output uart0_txd_o,
   output uart0_rts_o,
   output uart1_txd_o,
   output uart1_rts_o,
   output spi_clk_o,
   output spi_dat_o,
   output [7:0] spi_csn_o,
   output sdi_dat_o,
   output twi_sda_o,
   output twi_scl_o,
   output onewire_o,
   output [11:0] pwm_o,
   output [31:0] cfs_out_o,
   output neoled_o);
  wire [3:0] rstn_int_sreg;
  wire rstn_int;
  wire rstn_wdt;
  wire [11:0] clk_div;
  wire [11:0] clk_div_ff;
  wire [7:0] clk_gen;
  wire [10:0] clk_gen_en;
  wire clk_gen_en_ff;
  wire wdt_cg_en;
  wire uart0_cg_en;
  wire uart1_cg_en;
  wire spi_cg_en;
  wire twi_cg_en;
  wire pwm_cg_en;
  wire cfs_cg_en;
  wire neoled_cg_en;
  wire gptmr_cg_en;
  wire xip_cg_en;
  wire onewire_cg_en;
  wire [70:0] cpu_i;
  wire [70:0] i_cache;
  wire [107:0] cpu_d;
  wire [107:0] d_cache;
  wire [107:0] p_bus;
  wire bus_error;
  wire dci_ndmrstn;
  wire dci_halt_req;
  wire io_acc;
  wire io_rden;
  wire io_wren;
  reg [815:0] resp_bus;
  wire [15:0] fast_irq;
  wire mtime_irq;
  wire wdt_irq;
  wire uart0_rx_irq;
  wire uart0_tx_irq;
  wire uart1_rx_irq;
  wire uart1_tx_irq;
  wire spi_irq;
  wire sdi_irq;
  wire twi_irq;
  wire cfs_irq;
  wire neoled_irq;
  wire xirq_irq;
  wire gptmr_irq;
  wire onewire_irq;
  wire ext_timeout;
  wire ext_access;
  wire xip_access;
  wire xip_enable;
  wire [3:0] xip_page;
  wire n145_o;
  wire n150_o;
  wire n151_o;
  wire n152_o;
  wire [2:0] n153_o;
  wire [3:0] n155_o;
  wire [3:0] n157_o;
  wire n180_o;
  wire n182_o;
  wire n184_o;
  wire n185_o;
  wire n186_o;
  wire n187_o;
  wire n188_o;
  wire n189_o;
  wire n204_o;
  wire n212_o;
  wire n214_o;
  wire n216_o;
  wire n217_o;
  wire n218_o;
  wire n219_o;
  wire n220_o;
  wire n221_o;
  wire n222_o;
  wire n223_o;
  wire n224_o;
  wire n225_o;
  wire n226_o;
  wire n227_o;
  wire n228_o;
  wire n229_o;
  wire n230_o;
  wire n231_o;
  wire n232_o;
  wire n233_o;
  wire n234_o;
  wire n235_o;
  wire [11:0] n237_o;
  wire [11:0] n239_o;
  wire n250_o;
  wire n251_o;
  wire n252_o;
  wire n253_o;
  wire n254_o;
  wire n255_o;
  wire n256_o;
  wire n257_o;
  wire n258_o;
  wire n259_o;
  wire n260_o;
  wire n261_o;
  wire n262_o;
  wire n263_o;
  wire n264_o;
  wire n265_o;
  wire n266_o;
  wire n267_o;
  wire n268_o;
  wire n269_o;
  wire n270_o;
  wire n271_o;
  wire n272_o;
  wire n273_o;
  wire n274_o;
  wire n275_o;
  wire n276_o;
  wire n277_o;
  wire n278_o;
  wire n279_o;
  wire n280_o;
  wire n281_o;
  wire [31:0] neorv32_cpu_inst_n284;
  wire [31:0] n285_o;
  wire neorv32_cpu_inst_n286;
  wire n287_o;
  wire n288_o;
  wire neorv32_cpu_inst_n289;
  wire neorv32_cpu_inst_n290;
  wire [31:0] neorv32_cpu_inst_n291;
  wire [31:0] n292_o;
  wire [31:0] neorv32_cpu_inst_n293;
  wire [3:0] neorv32_cpu_inst_n294;
  wire neorv32_cpu_inst_n295;
  wire neorv32_cpu_inst_n296;
  wire n297_o;
  wire n298_o;
  wire neorv32_cpu_inst_n299;
  wire neorv32_cpu_inst_n300;
  wire neorv32_cpu_inst_sleep_o;
  wire neorv32_cpu_inst_debug_o;
  wire [31:0] neorv32_cpu_inst_i_bus_addr_o;
  wire neorv32_cpu_inst_i_bus_re_o;
  wire neorv32_cpu_inst_i_bus_fence_o;
  wire neorv32_cpu_inst_i_bus_priv_o;
  wire [31:0] neorv32_cpu_inst_d_bus_addr_o;
  wire [31:0] neorv32_cpu_inst_d_bus_wdata_o;
  wire [3:0] neorv32_cpu_inst_d_bus_ben_o;
  wire neorv32_cpu_inst_d_bus_we_o;
  wire neorv32_cpu_inst_d_bus_re_o;
  wire neorv32_cpu_inst_d_bus_fence_o;
  wire neorv32_cpu_inst_d_bus_priv_o;
  wire n331_o;
  wire n332_o;
  wire [31:0] n337_o;
  wire [31:0] n338_o;
  wire n339_o;
  wire n340_o;
  wire n341_o;
  wire n342_o;
  wire [31:0] n346_o;
  wire [31:0] n347_o;
  wire [31:0] n348_o;
  wire [3:0] n349_o;
  wire n350_o;
  wire n351_o;
  wire n352_o;
  wire n353_o;
  wire n354_o;
  wire n357_o;
  wire n358_o;
  wire [31:0] n359_o;
  wire [31:0] neorv32_busswitch_inst_n360;
  wire [31:0] n361_o;
  wire [3:0] n362_o;
  wire n363_o;
  wire n364_o;
  wire neorv32_busswitch_inst_n365;
  wire neorv32_busswitch_inst_n366;
  wire n367_o;
  wire n368_o;
  wire [31:0] n369_o;
  wire [31:0] neorv32_busswitch_inst_n370;
  localparam [31:0] n371_o = 32'b00000000000000000000000000000000;
  localparam [3:0] n372_o = 4'b0000;
  localparam n373_o = 1'b0;
  wire n374_o;
  wire neorv32_busswitch_inst_n375;
  wire neorv32_busswitch_inst_n376;
  wire neorv32_busswitch_inst_n377;
  wire neorv32_busswitch_inst_n378;
  wire neorv32_busswitch_inst_n379;
  wire [31:0] neorv32_busswitch_inst_n380;
  wire [31:0] n381_o;
  wire [31:0] neorv32_busswitch_inst_n382;
  wire [3:0] neorv32_busswitch_inst_n383;
  wire neorv32_busswitch_inst_n384;
  wire neorv32_busswitch_inst_n385;
  wire n386_o;
  wire [31:0] neorv32_busswitch_inst_ca_bus_rdata_o;
  wire neorv32_busswitch_inst_ca_bus_ack_o;
  wire neorv32_busswitch_inst_ca_bus_err_o;
  wire [31:0] neorv32_busswitch_inst_cb_bus_rdata_o;
  wire neorv32_busswitch_inst_cb_bus_ack_o;
  wire neorv32_busswitch_inst_cb_bus_err_o;
  wire neorv32_busswitch_inst_p_bus_priv_o;
  wire neorv32_busswitch_inst_p_bus_cached_o;
  wire neorv32_busswitch_inst_p_bus_src_o;
  wire [31:0] neorv32_busswitch_inst_p_bus_addr_o;
  wire [31:0] neorv32_busswitch_inst_p_bus_wdata_o;
  wire [3:0] neorv32_busswitch_inst_p_bus_ben_o;
  wire neorv32_busswitch_inst_p_bus_we_o;
  wire neorv32_busswitch_inst_p_bus_re_o;
  wire n415_o;
  wire n416_o;
  wire n417_o;
  wire [33:0] n422_o;
  wire [31:0] n423_o;
  wire [31:0] n425_o;
  wire [33:0] n427_o;
  wire n428_o;
  wire n430_o;
  wire [33:0] n432_o;
  wire n433_o;
  wire n435_o;
  wire [33:0] n437_o;
  wire [31:0] n438_o;
  wire [31:0] n439_o;
  wire [33:0] n440_o;
  wire n441_o;
  wire n442_o;
  wire [33:0] n443_o;
  wire n444_o;
  wire n445_o;
  wire [33:0] n446_o;
  wire [31:0] n447_o;
  wire [31:0] n448_o;
  wire [33:0] n449_o;
  wire n450_o;
  wire n451_o;
  wire [33:0] n452_o;
  wire n453_o;
  wire n454_o;
  wire [33:0] n455_o;
  wire [31:0] n456_o;
  wire [31:0] n457_o;
  wire [33:0] n458_o;
  wire n459_o;
  wire n460_o;
  wire [33:0] n461_o;
  wire n462_o;
  wire n463_o;
  wire [33:0] n464_o;
  wire [31:0] n465_o;
  wire [31:0] n466_o;
  wire [33:0] n467_o;
  wire n468_o;
  wire n469_o;
  wire [33:0] n470_o;
  wire n471_o;
  wire n472_o;
  wire [33:0] n473_o;
  wire [31:0] n474_o;
  wire [31:0] n475_o;
  wire [33:0] n476_o;
  wire n477_o;
  wire n478_o;
  wire [33:0] n479_o;
  wire n480_o;
  wire n481_o;
  wire [33:0] n482_o;
  wire [31:0] n483_o;
  wire [31:0] n484_o;
  wire [33:0] n485_o;
  wire n486_o;
  wire n487_o;
  wire [33:0] n488_o;
  wire n489_o;
  wire n490_o;
  wire [33:0] n491_o;
  wire [31:0] n492_o;
  wire [31:0] n493_o;
  wire [33:0] n494_o;
  wire n495_o;
  wire n496_o;
  wire [33:0] n497_o;
  wire n498_o;
  wire n499_o;
  wire [33:0] n500_o;
  wire [31:0] n501_o;
  wire [31:0] n502_o;
  wire [33:0] n503_o;
  wire n504_o;
  wire n505_o;
  wire [33:0] n506_o;
  wire n507_o;
  wire n508_o;
  wire [33:0] n509_o;
  wire [31:0] n510_o;
  wire [31:0] n511_o;
  wire [33:0] n512_o;
  wire n513_o;
  wire n514_o;
  wire [33:0] n515_o;
  wire n516_o;
  wire n517_o;
  wire [33:0] n518_o;
  wire [31:0] n519_o;
  wire [31:0] n520_o;
  wire [33:0] n521_o;
  wire n522_o;
  wire n523_o;
  wire [33:0] n524_o;
  wire n525_o;
  wire n526_o;
  wire [33:0] n527_o;
  wire [31:0] n528_o;
  wire [31:0] n529_o;
  wire [33:0] n530_o;
  wire n531_o;
  wire n532_o;
  wire [33:0] n533_o;
  wire n534_o;
  wire n535_o;
  wire [33:0] n536_o;
  wire [31:0] n537_o;
  wire [31:0] n538_o;
  wire [33:0] n539_o;
  wire n540_o;
  wire n541_o;
  wire [33:0] n542_o;
  wire n543_o;
  wire n544_o;
  wire [33:0] n545_o;
  wire [31:0] n546_o;
  wire [31:0] n547_o;
  wire [33:0] n548_o;
  wire n549_o;
  wire n550_o;
  wire [33:0] n551_o;
  wire n552_o;
  wire n553_o;
  wire [33:0] n554_o;
  wire [31:0] n555_o;
  wire [31:0] n556_o;
  wire [33:0] n557_o;
  wire n558_o;
  wire n559_o;
  wire [33:0] n560_o;
  wire n561_o;
  wire n562_o;
  wire [33:0] n563_o;
  wire [31:0] n564_o;
  wire [31:0] n565_o;
  wire [33:0] n566_o;
  wire n567_o;
  wire n568_o;
  wire [33:0] n569_o;
  wire n570_o;
  wire n571_o;
  wire [33:0] n572_o;
  wire [31:0] n573_o;
  wire [31:0] n574_o;
  wire [33:0] n575_o;
  wire n576_o;
  wire n577_o;
  wire [33:0] n578_o;
  wire n579_o;
  wire n580_o;
  wire [33:0] n581_o;
  wire [31:0] n582_o;
  wire [31:0] n583_o;
  wire [33:0] n584_o;
  wire n585_o;
  wire n586_o;
  wire [33:0] n587_o;
  wire n588_o;
  wire n589_o;
  wire [33:0] n590_o;
  wire [31:0] n591_o;
  wire [31:0] n592_o;
  wire [33:0] n593_o;
  wire n594_o;
  wire n595_o;
  wire [33:0] n596_o;
  wire n597_o;
  wire n598_o;
  wire [33:0] n599_o;
  wire [31:0] n600_o;
  wire [31:0] n601_o;
  wire [33:0] n602_o;
  wire n603_o;
  wire n604_o;
  wire [33:0] n605_o;
  wire n606_o;
  wire n607_o;
  wire [33:0] n608_o;
  wire [31:0] n609_o;
  wire [31:0] n610_o;
  wire [33:0] n611_o;
  wire n612_o;
  wire n613_o;
  wire [33:0] n614_o;
  wire n615_o;
  wire n616_o;
  wire [33:0] n617_o;
  wire [31:0] n618_o;
  wire [31:0] n619_o;
  wire [33:0] n620_o;
  wire n621_o;
  wire n622_o;
  wire [33:0] n623_o;
  wire n624_o;
  wire n625_o;
  wire [33:0] n626_o;
  wire [31:0] n627_o;
  wire [31:0] n628_o;
  wire [33:0] n629_o;
  wire n630_o;
  wire n631_o;
  wire [33:0] n632_o;
  wire n633_o;
  wire n634_o;
  wire [33:0] n635_o;
  wire [31:0] n636_o;
  wire [31:0] n637_o;
  wire [33:0] n638_o;
  wire n639_o;
  wire n640_o;
  wire [33:0] n641_o;
  wire n642_o;
  wire n643_o;
  wire [31:0] n645_o;
  wire [31:0] n646_o;
  wire [31:0] neorv32_bus_keeper_inst_n647;
  wire neorv32_bus_keeper_inst_n648;
  wire neorv32_bus_keeper_inst_n649;
  wire [31:0] n650_o;
  wire n651_o;
  wire n652_o;
  wire n653_o;
  wire n654_o;
  wire [31:0] neorv32_bus_keeper_inst_data_o;
  wire neorv32_bus_keeper_inst_ack_o;
  wire neorv32_bus_keeper_inst_err_o;
  wire n662_o;
  wire n663_o;
  wire [3:0] n664_o;
  wire [31:0] n665_o;
  wire [31:0] n666_o;
  wire [31:0] neorv32_int_imem_inst_true_neorv32_int_imem_inst_n667;
  wire neorv32_int_imem_inst_true_neorv32_int_imem_inst_n668;
  wire neorv32_int_imem_inst_true_neorv32_int_imem_inst_n669;
  wire [31:0] neorv32_int_imem_inst_true_neorv32_int_imem_inst_data_o;
  wire neorv32_int_imem_inst_true_neorv32_int_imem_inst_ack_o;
  wire neorv32_int_imem_inst_true_neorv32_int_imem_inst_err_o;
  wire n676_o;
  wire n677_o;
  wire [3:0] n678_o;
  wire [31:0] n679_o;
  wire [31:0] n680_o;
  wire [31:0] neorv32_int_dmem_inst_true_neorv32_int_dmem_inst_n681;
  wire neorv32_int_dmem_inst_true_neorv32_int_dmem_inst_n682;
  wire [31:0] neorv32_int_dmem_inst_true_neorv32_int_dmem_inst_data_o;
  wire neorv32_int_dmem_inst_true_neorv32_int_dmem_inst_ack_o;
  wire n688_o;
  wire n689_o;
  wire [31:0] n690_o;
  wire [31:0] neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_n691;
  wire neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_n692;
  wire neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_n693;
  wire [31:0] neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_data_o;
  wire neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_ack_o;
  wire neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_err_o;
  wire n700_o;
  wire [31:0] n701_o;
  wire n702_o;
  wire n703_o;
  wire [3:0] n704_o;
  wire [31:0] n705_o;
  wire [31:0] neorv32_wishbone_inst_true_neorv32_wishbone_inst_n706;
  wire neorv32_wishbone_inst_true_neorv32_wishbone_inst_n707;
  wire neorv32_wishbone_inst_true_neorv32_wishbone_inst_n708;
  wire neorv32_wishbone_inst_true_neorv32_wishbone_inst_n709;
  wire n710_o;
  wire neorv32_wishbone_inst_true_neorv32_wishbone_inst_n711;
  wire [2:0] neorv32_wishbone_inst_true_neorv32_wishbone_inst_n712;
  wire [31:0] neorv32_wishbone_inst_true_neorv32_wishbone_inst_n713;
  wire [31:0] neorv32_wishbone_inst_true_neorv32_wishbone_inst_n714;
  wire neorv32_wishbone_inst_true_neorv32_wishbone_inst_n715;
  wire [3:0] neorv32_wishbone_inst_true_neorv32_wishbone_inst_n716;
  wire neorv32_wishbone_inst_true_neorv32_wishbone_inst_n717;
  wire neorv32_wishbone_inst_true_neorv32_wishbone_inst_n718;
  wire [31:0] neorv32_wishbone_inst_true_neorv32_wishbone_inst_data_o;
  wire neorv32_wishbone_inst_true_neorv32_wishbone_inst_ack_o;
  wire neorv32_wishbone_inst_true_neorv32_wishbone_inst_err_o;
  wire neorv32_wishbone_inst_true_neorv32_wishbone_inst_tmo_o;
  wire neorv32_wishbone_inst_true_neorv32_wishbone_inst_ext_o;
  wire [2:0] neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_tag_o;
  wire [31:0] neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_adr_o;
  wire [31:0] neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_dat_o;
  wire neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_we_o;
  wire [3:0] neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_sel_o;
  wire neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_stb_o;
  wire neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_cyc_o;
  localparam n748_o = 1'b1;
  localparam n749_o = 1'b0;
  localparam n750_o = 1'b0;
  wire [22:0] n753_o;
  wire n756_o;
  wire n757_o;
  wire n760_o;
  wire n761_o;
  wire n762_o;
  wire n763_o;
  wire n764_o;
  wire n765_o;
  wire n768_o;
  wire n769_o;
  wire [3:0] n770_o;
  wire n772_o;
  wire n773_o;
  wire n774_o;
  localparam [31:0] n778_o = 32'b00000000000000000000000000000000;
  localparam n779_o = 1'b0;
  localparam [63:0] n781_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  wire [31:0] n785_o;
  wire [31:0] n786_o;
  wire [31:0] neorv32_mtime_inst_true_neorv32_mtime_inst_n787;
  wire neorv32_mtime_inst_true_neorv32_mtime_inst_n788;
  wire neorv32_mtime_inst_true_neorv32_mtime_inst_n789;
  wire [31:0] neorv32_mtime_inst_true_neorv32_mtime_inst_data_o;
  wire neorv32_mtime_inst_true_neorv32_mtime_inst_ack_o;
  wire neorv32_mtime_inst_true_neorv32_mtime_inst_irq_o;
  wire [31:0] n797_o;
  wire [31:0] n798_o;
  wire [31:0] neorv32_uart0_inst_true_neorv32_uart0_inst_n799;
  wire neorv32_uart0_inst_true_neorv32_uart0_inst_n800;
  wire neorv32_uart0_inst_true_neorv32_uart0_inst_n801;
  wire neorv32_uart0_inst_true_neorv32_uart0_inst_n802;
  wire neorv32_uart0_inst_true_neorv32_uart0_inst_n803;
  wire neorv32_uart0_inst_true_neorv32_uart0_inst_n804;
  wire neorv32_uart0_inst_true_neorv32_uart0_inst_n805;
  wire [31:0] neorv32_uart0_inst_true_neorv32_uart0_inst_data_o;
  wire neorv32_uart0_inst_true_neorv32_uart0_inst_ack_o;
  wire neorv32_uart0_inst_true_neorv32_uart0_inst_clkgen_en_o;
  wire neorv32_uart0_inst_true_neorv32_uart0_inst_uart_txd_o;
  wire neorv32_uart0_inst_true_neorv32_uart0_inst_uart_rts_o;
  wire neorv32_uart0_inst_true_neorv32_uart0_inst_irq_rx_o;
  wire neorv32_uart0_inst_true_neorv32_uart0_inst_irq_tx_o;
  localparam n821_o = 1'b0;
  localparam n822_o = 1'b1;
  localparam n826_o = 1'b0;
  localparam n827_o = 1'b0;
  localparam [7:0] n828_o = 8'b11111111;
  localparam n831_o = 1'b1;
  localparam n832_o = 1'b1;
  localparam [11:0] n836_o = 12'b000000000000;
  localparam n839_o = 1'b0;
  localparam n843_o = 1'b1;
  wire [31:0] n846_o;
  wire [31:0] neorv32_sysinfo_inst_n847;
  wire neorv32_sysinfo_inst_n848;
  wire neorv32_sysinfo_inst_n849;
  wire [31:0] neorv32_sysinfo_inst_data_o;
  wire neorv32_sysinfo_inst_ack_o;
  wire neorv32_sysinfo_inst_err_o;
  reg [3:0] n859_q;
  reg n861_q;
  reg [11:0] n862_q;
  reg [11:0] n863_q;
  wire [7:0] n864_o;
  wire [10:0] n865_o;
  reg n866_q;
  wire [70:0] n868_o;
  wire [70:0] n869_o;
  wire [107:0] n870_o;
  wire [107:0] n871_o;
  wire [107:0] n872_o;
  wire [815:0] n874_o;
  wire [15:0] n875_o;
  assign jtag_tdo_o = jtag_tdi_i;
  assign wb_tag_o = neorv32_wishbone_inst_true_neorv32_wishbone_inst_n712;
  assign wb_adr_o = neorv32_wishbone_inst_true_neorv32_wishbone_inst_n713;
  assign wb_dat_o = neorv32_wishbone_inst_true_neorv32_wishbone_inst_n714;
  assign wb_we_o = neorv32_wishbone_inst_true_neorv32_wishbone_inst_n715;
  assign wb_sel_o = neorv32_wishbone_inst_true_neorv32_wishbone_inst_n716;
  assign wb_stb_o = neorv32_wishbone_inst_true_neorv32_wishbone_inst_n717;
  assign wb_cyc_o = neorv32_wishbone_inst_true_neorv32_wishbone_inst_n718;
  assign fence_o = n331_o;
  assign fencei_o = n332_o;
  assign xip_csn_o = n748_o;
  assign xip_clk_o = n749_o;
  assign xip_dat_o = n750_o;
  assign gpio_o = n781_o;
  assign uart0_txd_o = neorv32_uart0_inst_true_neorv32_uart0_inst_n802;
  assign uart0_rts_o = neorv32_uart0_inst_true_neorv32_uart0_inst_n803;
  assign uart1_txd_o = n821_o;
  assign uart1_rts_o = n822_o;
  assign spi_clk_o = n826_o;
  assign spi_dat_o = n827_o;
  assign spi_csn_o = n828_o;
  assign sdi_dat_o = n779_o;
  assign twi_sda_o = n831_o;
  assign twi_scl_o = n832_o;
  assign onewire_o = n843_o;
  assign pwm_o = n836_o;
  assign cfs_out_o = n778_o;
  assign neoled_o = n839_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:245:10  */
  assign rstn_int_sreg = n859_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:247:10  */
  assign rstn_int = n861_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:248:10  */
  assign rstn_wdt = 1'b1; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:251:10  */
  assign clk_div = n862_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:252:10  */
  assign clk_div_ff = n863_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:253:10  */
  assign clk_gen = n864_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:254:10  */
  assign clk_gen_en = n865_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:255:10  */
  assign clk_gen_en_ff = n866_q; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:257:10  */
  assign wdt_cg_en = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:258:10  */
  assign uart0_cg_en = neorv32_uart0_inst_true_neorv32_uart0_inst_n801; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:259:10  */
  assign uart1_cg_en = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:260:10  */
  assign spi_cg_en = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:261:10  */
  assign twi_cg_en = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:262:10  */
  assign pwm_cg_en = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:263:10  */
  assign cfs_cg_en = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:264:10  */
  assign neoled_cg_en = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:265:10  */
  assign gptmr_cg_en = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:266:10  */
  assign xip_cg_en = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:267:10  */
  assign onewire_cg_en = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:288:10  */
  assign cpu_i = n868_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:288:17  */
  assign i_cache = n869_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:305:10  */
  assign cpu_d = n870_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:305:17  */
  assign d_cache = n871_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:305:26  */
  assign p_bus = n872_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:308:10  */
  assign bus_error = neorv32_bus_keeper_inst_n649; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:311:10  */
  assign dci_ndmrstn = 1'b1; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:312:10  */
  assign dci_halt_req = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:329:10  */
  assign io_acc = n757_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:330:10  */
  assign io_rden = n765_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:331:10  */
  assign io_wren = n774_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:351:10  */
  always @*
    resp_bus = n874_o; // (isignal)
  initial
    resp_bus = 816'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* ../neorv32/rtl/core/neorv32_top.vhd:354:10  */
  assign fast_irq = n875_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:355:10  */
  assign mtime_irq = neorv32_mtime_inst_true_neorv32_mtime_inst_n789; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:356:10  */
  assign wdt_irq = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:357:10  */
  assign uart0_rx_irq = neorv32_uart0_inst_true_neorv32_uart0_inst_n804; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:358:10  */
  assign uart0_tx_irq = neorv32_uart0_inst_true_neorv32_uart0_inst_n805; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:359:10  */
  assign uart1_rx_irq = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:360:10  */
  assign uart1_tx_irq = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:361:10  */
  assign spi_irq = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:362:10  */
  assign sdi_irq = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:363:10  */
  assign twi_irq = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:364:10  */
  assign cfs_irq = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:365:10  */
  assign neoled_irq = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:366:10  */
  assign xirq_irq = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:367:10  */
  assign gptmr_irq = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:368:10  */
  assign onewire_irq = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:371:10  */
  assign ext_timeout = neorv32_wishbone_inst_true_neorv32_wishbone_inst_n709; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:372:10  */
  assign ext_access = neorv32_wishbone_inst_true_neorv32_wishbone_inst_n711; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:373:10  */
  assign xip_access = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:374:10  */
  assign xip_enable = 1'b0; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:375:10  */
  assign xip_page = 4'b0000; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:444:16  */
  assign n145_o = ~rstn_i;
  /* ../neorv32/rtl/core/neorv32_top.vhd:453:20  */
  assign n150_o = ~rstn_wdt;
  /* ../neorv32/rtl/core/neorv32_top.vhd:453:43  */
  assign n151_o = ~dci_ndmrstn;
  /* ../neorv32/rtl/core/neorv32_top.vhd:453:27  */
  assign n152_o = n150_o | n151_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:456:39  */
  assign n153_o = rstn_int_sreg[2:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:456:71  */
  assign n155_o = {n153_o, 1'b1};
  /* ../neorv32/rtl/core/neorv32_top.vhd:453:7  */
  assign n157_o = n152_o ? 4'b0000 : n155_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2454:27  */
  assign n180_o = rstn_int_sreg[3];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2454:22  */
  assign n182_o = 1'b1 & n180_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2454:27  */
  assign n184_o = rstn_int_sreg[2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2454:22  */
  assign n185_o = n182_o & n184_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2454:27  */
  assign n186_o = rstn_int_sreg[1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2454:22  */
  assign n187_o = n185_o & n186_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2454:27  */
  assign n188_o = rstn_int_sreg[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2454:22  */
  assign n189_o = n187_o & n188_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:469:18  */
  assign n204_o = ~rstn_int;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n212_o = clk_gen_en[10];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n214_o = 1'b0 | n212_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n216_o = clk_gen_en[9];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n217_o = n214_o | n216_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n218_o = clk_gen_en[8];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n219_o = n217_o | n218_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n220_o = clk_gen_en[7];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n221_o = n219_o | n220_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n222_o = clk_gen_en[6];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n223_o = n221_o | n222_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n224_o = clk_gen_en[5];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n225_o = n223_o | n224_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n226_o = clk_gen_en[4];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n227_o = n225_o | n226_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n228_o = clk_gen_en[3];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n229_o = n227_o | n228_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n230_o = clk_gen_en[2];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n231_o = n229_o | n230_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n232_o = clk_gen_en[1];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n233_o = n231_o | n232_o;
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:26  */
  assign n234_o = clk_gen_en[0];
  /* ../neorv32/rtl/core/neorv32_package.vhd:2442:22  */
  assign n235_o = n233_o | n234_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:476:56  */
  assign n237_o = clk_div + 12'b000000000001;
  /* ../neorv32/rtl/core/neorv32_top.vhd:475:7  */
  assign n239_o = clk_gen_en_ff ? n237_o : 12'b000000000000;
  /* ../neorv32/rtl/core/neorv32_top.vhd:485:36  */
  assign n250_o = clk_div[0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:485:60  */
  assign n251_o = clk_div_ff[0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:485:46  */
  assign n252_o = ~n251_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:485:41  */
  assign n253_o = n250_o & n252_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:486:36  */
  assign n254_o = clk_div[1];
  /* ../neorv32/rtl/core/neorv32_top.vhd:486:60  */
  assign n255_o = clk_div_ff[1];
  /* ../neorv32/rtl/core/neorv32_top.vhd:486:46  */
  assign n256_o = ~n255_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:486:41  */
  assign n257_o = n254_o & n256_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:487:36  */
  assign n258_o = clk_div[2];
  /* ../neorv32/rtl/core/neorv32_top.vhd:487:60  */
  assign n259_o = clk_div_ff[2];
  /* ../neorv32/rtl/core/neorv32_top.vhd:487:46  */
  assign n260_o = ~n259_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:487:41  */
  assign n261_o = n258_o & n260_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:488:36  */
  assign n262_o = clk_div[5];
  /* ../neorv32/rtl/core/neorv32_top.vhd:488:60  */
  assign n263_o = clk_div_ff[5];
  /* ../neorv32/rtl/core/neorv32_top.vhd:488:46  */
  assign n264_o = ~n263_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:488:41  */
  assign n265_o = n262_o & n264_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:489:36  */
  assign n266_o = clk_div[6];
  /* ../neorv32/rtl/core/neorv32_top.vhd:489:60  */
  assign n267_o = clk_div_ff[6];
  /* ../neorv32/rtl/core/neorv32_top.vhd:489:46  */
  assign n268_o = ~n267_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:489:41  */
  assign n269_o = n266_o & n268_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:490:36  */
  assign n270_o = clk_div[9];
  /* ../neorv32/rtl/core/neorv32_top.vhd:490:60  */
  assign n271_o = clk_div_ff[9];
  /* ../neorv32/rtl/core/neorv32_top.vhd:490:46  */
  assign n272_o = ~n271_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:490:41  */
  assign n273_o = n270_o & n272_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:491:36  */
  assign n274_o = clk_div[10];
  /* ../neorv32/rtl/core/neorv32_top.vhd:491:60  */
  assign n275_o = clk_div_ff[10];
  /* ../neorv32/rtl/core/neorv32_top.vhd:491:46  */
  assign n276_o = ~n275_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:491:41  */
  assign n277_o = n274_o & n276_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:492:36  */
  assign n278_o = clk_div[11];
  /* ../neorv32/rtl/core/neorv32_top.vhd:492:60  */
  assign n279_o = clk_div_ff[11];
  /* ../neorv32/rtl/core/neorv32_top.vhd:492:46  */
  assign n280_o = ~n279_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:492:41  */
  assign n281_o = n278_o & n280_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:555:22  */
  assign neorv32_cpu_inst_n284 = neorv32_cpu_inst_i_bus_addr_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:556:28  */
  assign n285_o = cpu_i[63:32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:557:22  */
  assign neorv32_cpu_inst_n286 = neorv32_cpu_inst_i_bus_re_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:558:28  */
  assign n287_o = cpu_i[65];
  /* ../neorv32/rtl/core/neorv32_top.vhd:559:28  */
  assign n288_o = cpu_i[66];
  /* ../neorv32/rtl/core/neorv32_top.vhd:560:22  */
  assign neorv32_cpu_inst_n289 = neorv32_cpu_inst_i_bus_fence_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:561:22  */
  assign neorv32_cpu_inst_n290 = neorv32_cpu_inst_i_bus_priv_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:563:22  */
  assign neorv32_cpu_inst_n291 = neorv32_cpu_inst_d_bus_addr_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:564:28  */
  assign n292_o = cpu_d[63:32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:565:22  */
  assign neorv32_cpu_inst_n293 = neorv32_cpu_inst_d_bus_wdata_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:566:22  */
  assign neorv32_cpu_inst_n294 = neorv32_cpu_inst_d_bus_ben_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:567:22  */
  assign neorv32_cpu_inst_n295 = neorv32_cpu_inst_d_bus_we_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:568:22  */
  assign neorv32_cpu_inst_n296 = neorv32_cpu_inst_d_bus_re_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:569:28  */
  assign n297_o = cpu_d[102];
  /* ../neorv32/rtl/core/neorv32_top.vhd:570:28  */
  assign n298_o = cpu_d[103];
  /* ../neorv32/rtl/core/neorv32_top.vhd:571:22  */
  assign neorv32_cpu_inst_n299 = neorv32_cpu_inst_d_bus_fence_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:572:22  */
  assign neorv32_cpu_inst_n300 = neorv32_cpu_inst_d_bus_priv_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:514:3  */
  neorv32_cpu_1_0_4_0_40_8cd82fcc1d144656bad81224642c94d0248852b6 neorv32_cpu_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_int),
    .i_bus_rdata_i(n285_o),
    .i_bus_ack_i(n287_o),
    .i_bus_err_i(n288_o),
    .d_bus_rdata_i(n292_o),
    .d_bus_ack_i(n297_o),
    .d_bus_err_i(n298_o),
    .msw_irq_i(msw_irq_i),
    .mext_irq_i(mext_irq_i),
    .mtime_irq_i(mtime_irq),
    .firq_i(fast_irq),
    .db_halt_req_i(dci_halt_req),
    .sleep_o(),
    .debug_o(),
    .i_bus_addr_o(neorv32_cpu_inst_i_bus_addr_o),
    .i_bus_re_o(neorv32_cpu_inst_i_bus_re_o),
    .i_bus_fence_o(neorv32_cpu_inst_i_bus_fence_o),
    .i_bus_priv_o(neorv32_cpu_inst_i_bus_priv_o),
    .d_bus_addr_o(neorv32_cpu_inst_d_bus_addr_o),
    .d_bus_wdata_o(neorv32_cpu_inst_d_bus_wdata_o),
    .d_bus_ben_o(neorv32_cpu_inst_d_bus_ben_o),
    .d_bus_we_o(neorv32_cpu_inst_d_bus_we_o),
    .d_bus_re_o(neorv32_cpu_inst_d_bus_re_o),
    .d_bus_fence_o(neorv32_cpu_inst_d_bus_fence_o),
    .d_bus_priv_o(neorv32_cpu_inst_d_bus_priv_o));
  /* ../neorv32/rtl/core/neorv32_top.vhd:590:21  */
  assign n331_o = cpu_d[104];
  /* ../neorv32/rtl/core/neorv32_top.vhd:591:21  */
  assign n332_o = cpu_i[67];
  /* ../neorv32/rtl/core/neorv32_top.vhd:646:29  */
  assign n337_o = cpu_i[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:647:31  */
  assign n338_o = i_cache[63:32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:648:29  */
  assign n339_o = cpu_i[64];
  /* ../neorv32/rtl/core/neorv32_top.vhd:649:31  */
  assign n340_o = i_cache[65];
  /* ../neorv32/rtl/core/neorv32_top.vhd:650:31  */
  assign n341_o = i_cache[66];
  /* ../neorv32/rtl/core/neorv32_top.vhd:653:26  */
  assign n342_o = cpu_i[70];
  /* ../neorv32/rtl/core/neorv32_top.vhd:698:29  */
  assign n346_o = cpu_d[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:699:31  */
  assign n347_o = d_cache[63:32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:700:29  */
  assign n348_o = cpu_d[95:64];
  /* ../neorv32/rtl/core/neorv32_top.vhd:701:29  */
  assign n349_o = cpu_d[99:96];
  /* ../neorv32/rtl/core/neorv32_top.vhd:702:29  */
  assign n350_o = cpu_d[100];
  /* ../neorv32/rtl/core/neorv32_top.vhd:703:29  */
  assign n351_o = cpu_d[101];
  /* ../neorv32/rtl/core/neorv32_top.vhd:704:31  */
  assign n352_o = d_cache[102];
  /* ../neorv32/rtl/core/neorv32_top.vhd:705:31  */
  assign n353_o = d_cache[103];
  /* ../neorv32/rtl/core/neorv32_top.vhd:708:26  */
  assign n354_o = cpu_d[107];
  /* ../neorv32/rtl/core/neorv32_top.vhd:725:32  */
  assign n357_o = d_cache[107];
  /* ../neorv32/rtl/core/neorv32_top.vhd:726:32  */
  assign n358_o = d_cache[106];
  /* ../neorv32/rtl/core/neorv32_top.vhd:727:32  */
  assign n359_o = d_cache[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:728:24  */
  assign neorv32_busswitch_inst_n360 = neorv32_busswitch_inst_ca_bus_rdata_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:729:32  */
  assign n361_o = d_cache[95:64];
  /* ../neorv32/rtl/core/neorv32_top.vhd:730:32  */
  assign n362_o = d_cache[99:96];
  /* ../neorv32/rtl/core/neorv32_top.vhd:731:32  */
  assign n363_o = d_cache[100];
  /* ../neorv32/rtl/core/neorv32_top.vhd:732:32  */
  assign n364_o = d_cache[101];
  /* ../neorv32/rtl/core/neorv32_top.vhd:733:24  */
  assign neorv32_busswitch_inst_n365 = neorv32_busswitch_inst_ca_bus_ack_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:734:24  */
  assign neorv32_busswitch_inst_n366 = neorv32_busswitch_inst_ca_bus_err_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:736:32  */
  assign n367_o = i_cache[70];
  /* ../neorv32/rtl/core/neorv32_top.vhd:737:32  */
  assign n368_o = i_cache[69];
  /* ../neorv32/rtl/core/neorv32_top.vhd:738:32  */
  assign n369_o = i_cache[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:739:24  */
  assign neorv32_busswitch_inst_n370 = neorv32_busswitch_inst_cb_bus_rdata_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:743:32  */
  assign n374_o = i_cache[64];
  /* ../neorv32/rtl/core/neorv32_top.vhd:744:24  */
  assign neorv32_busswitch_inst_n375 = neorv32_busswitch_inst_cb_bus_ack_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:745:24  */
  assign neorv32_busswitch_inst_n376 = neorv32_busswitch_inst_cb_bus_err_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:747:24  */
  assign neorv32_busswitch_inst_n377 = neorv32_busswitch_inst_p_bus_priv_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:748:24  */
  assign neorv32_busswitch_inst_n378 = neorv32_busswitch_inst_p_bus_cached_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:749:24  */
  assign neorv32_busswitch_inst_n379 = neorv32_busswitch_inst_p_bus_src_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:750:24  */
  assign neorv32_busswitch_inst_n380 = neorv32_busswitch_inst_p_bus_addr_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:751:30  */
  assign n381_o = p_bus[63:32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:752:24  */
  assign neorv32_busswitch_inst_n382 = neorv32_busswitch_inst_p_bus_wdata_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:753:24  */
  assign neorv32_busswitch_inst_n383 = neorv32_busswitch_inst_p_bus_ben_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:754:24  */
  assign neorv32_busswitch_inst_n384 = neorv32_busswitch_inst_p_bus_we_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:755:24  */
  assign neorv32_busswitch_inst_n385 = neorv32_busswitch_inst_p_bus_re_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:756:30  */
  assign n386_o = p_bus[102];
  /* ../neorv32/rtl/core/neorv32_top.vhd:715:3  */
  neorv32_busswitch_3f29546453678b855931c174a97d6c0894b8f546 neorv32_busswitch_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_int),
    .ca_bus_priv_i(n357_o),
    .ca_bus_cached_i(n358_o),
    .ca_bus_addr_i(n359_o),
    .ca_bus_wdata_i(n361_o),
    .ca_bus_ben_i(n362_o),
    .ca_bus_we_i(n363_o),
    .ca_bus_re_i(n364_o),
    .cb_bus_priv_i(n367_o),
    .cb_bus_cached_i(n368_o),
    .cb_bus_addr_i(n369_o),
    .cb_bus_wdata_i(n371_o),
    .cb_bus_ben_i(n372_o),
    .cb_bus_we_i(n373_o),
    .cb_bus_re_i(n374_o),
    .p_bus_rdata_i(n381_o),
    .p_bus_ack_i(n386_o),
    .p_bus_err_i(bus_error),
    .ca_bus_rdata_o(neorv32_busswitch_inst_ca_bus_rdata_o),
    .ca_bus_ack_o(neorv32_busswitch_inst_ca_bus_ack_o),
    .ca_bus_err_o(neorv32_busswitch_inst_ca_bus_err_o),
    .cb_bus_rdata_o(neorv32_busswitch_inst_cb_bus_rdata_o),
    .cb_bus_ack_o(neorv32_busswitch_inst_cb_bus_ack_o),
    .cb_bus_err_o(neorv32_busswitch_inst_cb_bus_err_o),
    .p_bus_priv_o(neorv32_busswitch_inst_p_bus_priv_o),
    .p_bus_cached_o(neorv32_busswitch_inst_p_bus_cached_o),
    .p_bus_src_o(neorv32_busswitch_inst_p_bus_src_o),
    .p_bus_addr_o(neorv32_busswitch_inst_p_bus_addr_o),
    .p_bus_wdata_o(neorv32_busswitch_inst_p_bus_wdata_o),
    .p_bus_ben_o(neorv32_busswitch_inst_p_bus_ben_o),
    .p_bus_we_o(neorv32_busswitch_inst_p_bus_we_o),
    .p_bus_re_o(neorv32_busswitch_inst_p_bus_re_o));
  /* ../neorv32/rtl/core/neorv32_top.vhd:761:24  */
  assign n415_o = cpu_i[67];
  /* ../neorv32/rtl/core/neorv32_top.vhd:761:39  */
  assign n416_o = cpu_d[104];
  /* ../neorv32/rtl/core/neorv32_top.vhd:761:30  */
  assign n417_o = n415_o | n416_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n422_o = resp_bus[815:782];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n423_o = n422_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n425_o = 32'b00000000000000000000000000000000 | n423_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n427_o = resp_bus[815:782];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n428_o = n427_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n430_o = 1'b0 | n428_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n432_o = resp_bus[815:782];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n433_o = n432_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n435_o = 1'b0 | n433_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n437_o = resp_bus[781:748];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n438_o = n437_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n439_o = n425_o | n438_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n440_o = resp_bus[781:748];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n441_o = n440_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n442_o = n430_o | n441_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n443_o = resp_bus[781:748];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n444_o = n443_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n445_o = n435_o | n444_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n446_o = resp_bus[747:714];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n447_o = n446_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n448_o = n439_o | n447_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n449_o = resp_bus[747:714];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n450_o = n449_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n451_o = n442_o | n450_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n452_o = resp_bus[747:714];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n453_o = n452_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n454_o = n445_o | n453_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n455_o = resp_bus[713:680];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n456_o = n455_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n457_o = n448_o | n456_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n458_o = resp_bus[713:680];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n459_o = n458_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n460_o = n451_o | n459_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n461_o = resp_bus[713:680];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n462_o = n461_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n463_o = n454_o | n462_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n464_o = resp_bus[679:646];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n465_o = n464_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n466_o = n457_o | n465_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n467_o = resp_bus[679:646];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n468_o = n467_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n469_o = n460_o | n468_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n470_o = resp_bus[679:646];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n471_o = n470_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n472_o = n463_o | n471_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n473_o = resp_bus[645:612];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n474_o = n473_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n475_o = n466_o | n474_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n476_o = resp_bus[645:612];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n477_o = n476_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n478_o = n469_o | n477_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n479_o = resp_bus[645:612];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n480_o = n479_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n481_o = n472_o | n480_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n482_o = resp_bus[611:578];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n483_o = n482_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n484_o = n475_o | n483_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n485_o = resp_bus[611:578];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n486_o = n485_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n487_o = n478_o | n486_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n488_o = resp_bus[611:578];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n489_o = n488_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n490_o = n481_o | n489_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n491_o = resp_bus[577:544];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n492_o = n491_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n493_o = n484_o | n492_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n494_o = resp_bus[577:544];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n495_o = n494_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n496_o = n487_o | n495_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n497_o = resp_bus[577:544];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n498_o = n497_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n499_o = n490_o | n498_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n500_o = resp_bus[543:510];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n501_o = n500_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n502_o = n493_o | n501_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n503_o = resp_bus[543:510];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n504_o = n503_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n505_o = n496_o | n504_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n506_o = resp_bus[543:510];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n507_o = n506_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n508_o = n499_o | n507_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n509_o = resp_bus[509:476];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n510_o = n509_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n511_o = n502_o | n510_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n512_o = resp_bus[509:476];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n513_o = n512_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n514_o = n505_o | n513_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n515_o = resp_bus[509:476];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n516_o = n515_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n517_o = n508_o | n516_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n518_o = resp_bus[475:442];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n519_o = n518_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n520_o = n511_o | n519_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n521_o = resp_bus[475:442];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n522_o = n521_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n523_o = n514_o | n522_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n524_o = resp_bus[475:442];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n525_o = n524_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n526_o = n517_o | n525_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n527_o = resp_bus[441:408];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n528_o = n527_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n529_o = n520_o | n528_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n530_o = resp_bus[441:408];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n531_o = n530_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n532_o = n523_o | n531_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n533_o = resp_bus[441:408];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n534_o = n533_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n535_o = n526_o | n534_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n536_o = resp_bus[407:374];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n537_o = n536_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n538_o = n529_o | n537_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n539_o = resp_bus[407:374];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n540_o = n539_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n541_o = n532_o | n540_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n542_o = resp_bus[407:374];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n543_o = n542_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n544_o = n535_o | n543_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n545_o = resp_bus[373:340];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n546_o = n545_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n547_o = n538_o | n546_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n548_o = resp_bus[373:340];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n549_o = n548_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n550_o = n541_o | n549_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n551_o = resp_bus[373:340];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n552_o = n551_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n553_o = n544_o | n552_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n554_o = resp_bus[339:306];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n555_o = n554_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n556_o = n547_o | n555_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n557_o = resp_bus[339:306];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n558_o = n557_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n559_o = n550_o | n558_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n560_o = resp_bus[339:306];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n561_o = n560_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n562_o = n553_o | n561_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n563_o = resp_bus[305:272];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n564_o = n563_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n565_o = n556_o | n564_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n566_o = resp_bus[305:272];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n567_o = n566_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n568_o = n559_o | n567_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n569_o = resp_bus[305:272];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n570_o = n569_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n571_o = n562_o | n570_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n572_o = resp_bus[271:238];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n573_o = n572_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n574_o = n565_o | n573_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n575_o = resp_bus[271:238];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n576_o = n575_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n577_o = n568_o | n576_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n578_o = resp_bus[271:238];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n579_o = n578_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n580_o = n571_o | n579_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n581_o = resp_bus[237:204];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n582_o = n581_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n583_o = n574_o | n582_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n584_o = resp_bus[237:204];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n585_o = n584_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n586_o = n577_o | n585_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n587_o = resp_bus[237:204];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n588_o = n587_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n589_o = n580_o | n588_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n590_o = resp_bus[203:170];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n591_o = n590_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n592_o = n583_o | n591_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n593_o = resp_bus[203:170];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n594_o = n593_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n595_o = n586_o | n594_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n596_o = resp_bus[203:170];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n597_o = n596_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n598_o = n589_o | n597_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n599_o = resp_bus[169:136];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n600_o = n599_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n601_o = n592_o | n600_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n602_o = resp_bus[169:136];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n603_o = n602_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n604_o = n595_o | n603_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n605_o = resp_bus[169:136];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n606_o = n605_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n607_o = n598_o | n606_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n608_o = resp_bus[135:102];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n609_o = n608_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n610_o = n601_o | n609_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n611_o = resp_bus[135:102];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n612_o = n611_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n613_o = n604_o | n612_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n614_o = resp_bus[135:102];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n615_o = n614_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n616_o = n607_o | n615_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n617_o = resp_bus[101:68];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n618_o = n617_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n619_o = n610_o | n618_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n620_o = resp_bus[101:68];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n621_o = n620_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n622_o = n613_o | n621_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n623_o = resp_bus[101:68];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n624_o = n623_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n625_o = n616_o | n624_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n626_o = resp_bus[67:34];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n627_o = n626_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n628_o = n619_o | n627_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n629_o = resp_bus[67:34];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n630_o = n629_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n631_o = n622_o | n630_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n632_o = resp_bus[67:34];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n633_o = n632_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n634_o = n625_o | n633_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:37  */
  assign n635_o = resp_bus[33:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:41  */
  assign n636_o = n635_o[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:775:26  */
  assign n637_o = n628_o | n636_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:37  */
  assign n638_o = resp_bus[33:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:41  */
  assign n639_o = n638_o[32];
  /* ../neorv32/rtl/core/neorv32_top.vhd:776:26  */
  assign n640_o = n631_o | n639_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:37  */
  assign n641_o = resp_bus[33:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:41  */
  assign n642_o = n641_o[33];
  /* ../neorv32/rtl/core/neorv32_top.vhd:777:26  */
  assign n643_o = n634_o | n642_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:792:25  */
  assign n645_o = p_bus[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:795:25  */
  assign n646_o = p_bus[95:64];
  /* ../neorv32/rtl/core/neorv32_top.vhd:796:19  */
  assign neorv32_bus_keeper_inst_n647 = neorv32_bus_keeper_inst_data_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:797:19  */
  assign neorv32_bus_keeper_inst_n648 = neorv32_bus_keeper_inst_ack_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:798:19  */
  assign neorv32_bus_keeper_inst_n649 = neorv32_bus_keeper_inst_err_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:800:25  */
  assign n650_o = p_bus[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:801:25  */
  assign n651_o = p_bus[101];
  /* ../neorv32/rtl/core/neorv32_top.vhd:802:25  */
  assign n652_o = p_bus[100];
  /* ../neorv32/rtl/core/neorv32_top.vhd:803:25  */
  assign n653_o = p_bus[102];
  /* ../neorv32/rtl/core/neorv32_top.vhd:804:25  */
  assign n654_o = p_bus[103];
  /* ../neorv32/rtl/core/neorv32_top.vhd:787:3  */
  neorv32_bus_keeper neorv32_bus_keeper_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_int),
    .addr_i(n645_o),
    .rden_i(io_rden),
    .wren_i(io_wren),
    .data_i(n646_o),
    .bus_addr_i(n650_o),
    .bus_rden_i(n651_o),
    .bus_wren_i(n652_o),
    .bus_ack_i(n653_o),
    .bus_err_i(n654_o),
    .bus_tmo_i(ext_timeout),
    .bus_ext_i(ext_access),
    .bus_xip_i(xip_access),
    .data_o(neorv32_bus_keeper_inst_data_o),
    .ack_o(neorv32_bus_keeper_inst_ack_o),
    .err_o(neorv32_bus_keeper_inst_err_o));
  /* ../neorv32/rtl/core/neorv32_top.vhd:830:23  */
  assign n662_o = p_bus[101];
  /* ../neorv32/rtl/core/neorv32_top.vhd:831:23  */
  assign n663_o = p_bus[100];
  /* ../neorv32/rtl/core/neorv32_top.vhd:832:23  */
  assign n664_o = p_bus[99:96];
  /* ../neorv32/rtl/core/neorv32_top.vhd:833:23  */
  assign n665_o = p_bus[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:834:23  */
  assign n666_o = p_bus[95:64];
  /* ../neorv32/rtl/core/neorv32_top.vhd:835:17  */
  assign neorv32_int_imem_inst_true_neorv32_int_imem_inst_n667 = neorv32_int_imem_inst_true_neorv32_int_imem_inst_data_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:836:17  */
  assign neorv32_int_imem_inst_true_neorv32_int_imem_inst_n668 = neorv32_int_imem_inst_true_neorv32_int_imem_inst_ack_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:837:17  */
  assign neorv32_int_imem_inst_true_neorv32_int_imem_inst_n669 = neorv32_int_imem_inst_true_neorv32_int_imem_inst_err_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:822:5  */
  neorv32_imem_1024_91a7f356ca6ce41b6122bd41e60c1f2eb8f0f0e3 neorv32_int_imem_inst_true_neorv32_int_imem_inst (
    .clk_i(clk_i),
    .rden_i(n662_o),
    .wren_i(n663_o),
    .ben_i(n664_o),
    .addr_i(n665_o),
    .data_i(n666_o),
    .data_o(neorv32_int_imem_inst_true_neorv32_int_imem_inst_data_o),
    .ack_o(neorv32_int_imem_inst_true_neorv32_int_imem_inst_ack_o),
    .err_o(neorv32_int_imem_inst_true_neorv32_int_imem_inst_err_o));
  /* ../neorv32/rtl/core/neorv32_top.vhd:858:23  */
  assign n676_o = p_bus[101];
  /* ../neorv32/rtl/core/neorv32_top.vhd:859:23  */
  assign n677_o = p_bus[100];
  /* ../neorv32/rtl/core/neorv32_top.vhd:860:23  */
  assign n678_o = p_bus[99:96];
  /* ../neorv32/rtl/core/neorv32_top.vhd:861:23  */
  assign n679_o = p_bus[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:862:23  */
  assign n680_o = p_bus[95:64];
  /* ../neorv32/rtl/core/neorv32_top.vhd:863:17  */
  assign neorv32_int_dmem_inst_true_neorv32_int_dmem_inst_n681 = neorv32_int_dmem_inst_true_neorv32_int_dmem_inst_data_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:864:17  */
  assign neorv32_int_dmem_inst_true_neorv32_int_dmem_inst_n682 = neorv32_int_dmem_inst_true_neorv32_int_dmem_inst_ack_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:851:5  */
  neorv32_dmem_2048_34d7de1b571aa545cf571b84dc4b40d1f42fed39 neorv32_int_dmem_inst_true_neorv32_int_dmem_inst (
    .clk_i(clk_i),
    .rden_i(n676_o),
    .wren_i(n677_o),
    .ben_i(n678_o),
    .addr_i(n679_o),
    .data_i(n680_o),
    .data_o(neorv32_int_dmem_inst_true_neorv32_int_dmem_inst_data_o),
    .ack_o(neorv32_int_dmem_inst_true_neorv32_int_dmem_inst_ack_o));
  /* ../neorv32/rtl/core/neorv32_top.vhd:885:23  */
  assign n688_o = p_bus[101];
  /* ../neorv32/rtl/core/neorv32_top.vhd:886:23  */
  assign n689_o = p_bus[100];
  /* ../neorv32/rtl/core/neorv32_top.vhd:887:23  */
  assign n690_o = p_bus[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:888:17  */
  assign neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_n691 = neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_data_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:889:17  */
  assign neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_n692 = neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_ack_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:890:17  */
  assign neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_n693 = neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_err_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:879:5  */
  neorv32_boot_rom_8aaa057a3ce108fd664b4f820549d0c7a5c85d77 neorv32_boot_rom_inst_true_neorv32_boot_rom_inst (
    .clk_i(clk_i),
    .rden_i(n688_o),
    .wren_i(n689_o),
    .addr_i(n690_o),
    .data_o(neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_data_o),
    .ack_o(neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_ack_o),
    .err_o(neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_err_o));
  /* ../neorv32/rtl/core/neorv32_top.vhd:924:27  */
  assign n700_o = p_bus[105];
  /* ../neorv32/rtl/core/neorv32_top.vhd:925:27  */
  assign n701_o = p_bus[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:926:27  */
  assign n702_o = p_bus[101];
  /* ../neorv32/rtl/core/neorv32_top.vhd:927:27  */
  assign n703_o = p_bus[100];
  /* ../neorv32/rtl/core/neorv32_top.vhd:928:27  */
  assign n704_o = p_bus[99:96];
  /* ../neorv32/rtl/core/neorv32_top.vhd:929:27  */
  assign n705_o = p_bus[95:64];
  /* ../neorv32/rtl/core/neorv32_top.vhd:930:21  */
  assign neorv32_wishbone_inst_true_neorv32_wishbone_inst_n706 = neorv32_wishbone_inst_true_neorv32_wishbone_inst_data_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:931:21  */
  assign neorv32_wishbone_inst_true_neorv32_wishbone_inst_n707 = neorv32_wishbone_inst_true_neorv32_wishbone_inst_ack_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:932:21  */
  assign neorv32_wishbone_inst_true_neorv32_wishbone_inst_n708 = neorv32_wishbone_inst_true_neorv32_wishbone_inst_err_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:933:21  */
  assign neorv32_wishbone_inst_true_neorv32_wishbone_inst_n709 = neorv32_wishbone_inst_true_neorv32_wishbone_inst_tmo_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:934:27  */
  assign n710_o = p_bus[107];
  /* ../neorv32/rtl/core/neorv32_top.vhd:935:21  */
  assign neorv32_wishbone_inst_true_neorv32_wishbone_inst_n711 = neorv32_wishbone_inst_true_neorv32_wishbone_inst_ext_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:940:21  */
  assign neorv32_wishbone_inst_true_neorv32_wishbone_inst_n712 = neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_tag_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:941:21  */
  assign neorv32_wishbone_inst_true_neorv32_wishbone_inst_n713 = neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_adr_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:943:21  */
  assign neorv32_wishbone_inst_true_neorv32_wishbone_inst_n714 = neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_dat_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:944:21  */
  assign neorv32_wishbone_inst_true_neorv32_wishbone_inst_n715 = neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_we_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:945:21  */
  assign neorv32_wishbone_inst_true_neorv32_wishbone_inst_n716 = neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_sel_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:946:21  */
  assign neorv32_wishbone_inst_true_neorv32_wishbone_inst_n717 = neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_stb_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:947:21  */
  assign neorv32_wishbone_inst_true_neorv32_wishbone_inst_n718 = neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_cyc_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:904:5  */
  neorv32_wishbone_1024_2048_255_faf1cd4bdf2d59261beed066baf3c3e69ee5d9f7 neorv32_wishbone_inst_true_neorv32_wishbone_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_int),
    .src_i(n700_o),
    .addr_i(n701_o),
    .rden_i(n702_o),
    .wren_i(n703_o),
    .ben_i(n704_o),
    .data_i(n705_o),
    .priv_i(n710_o),
    .xip_en_i(xip_enable),
    .xip_page_i(xip_page),
    .wb_dat_i(wb_dat_i),
    .wb_ack_i(wb_ack_i),
    .wb_err_i(wb_err_i),
    .data_o(neorv32_wishbone_inst_true_neorv32_wishbone_inst_data_o),
    .ack_o(neorv32_wishbone_inst_true_neorv32_wishbone_inst_ack_o),
    .err_o(neorv32_wishbone_inst_true_neorv32_wishbone_inst_err_o),
    .tmo_o(neorv32_wishbone_inst_true_neorv32_wishbone_inst_tmo_o),
    .ext_o(neorv32_wishbone_inst_true_neorv32_wishbone_inst_ext_o),
    .wb_tag_o(neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_tag_o),
    .wb_adr_o(neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_adr_o),
    .wb_dat_o(neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_dat_o),
    .wb_we_o(neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_we_o),
    .wb_sel_o(neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_sel_o),
    .wb_stb_o(neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_stb_o),
    .wb_cyc_o(neorv32_wishbone_inst_true_neorv32_wishbone_inst_wb_cyc_o));
  /* ../neorv32/rtl/core/neorv32_top.vhd:1029:34  */
  assign n753_o = p_bus[31:9];
  /* ../neorv32/rtl/core/neorv32_top.vhd:1029:70  */
  assign n756_o = n753_o == 23'b11111111111111111111111;
  /* ../neorv32/rtl/core/neorv32_top.vhd:1029:18  */
  assign n757_o = n756_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_top.vhd:1030:49  */
  assign n760_o = p_bus[101];
  /* ../neorv32/rtl/core/neorv32_top.vhd:1030:38  */
  assign n761_o = io_acc & n760_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:1030:70  */
  assign n762_o = p_bus[105];
  /* ../neorv32/rtl/core/neorv32_top.vhd:1030:74  */
  assign n763_o = ~n762_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:1030:59  */
  assign n764_o = n761_o & n763_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:1030:18  */
  assign n765_o = n764_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_top.vhd:1031:49  */
  assign n768_o = p_bus[100];
  /* ../neorv32/rtl/core/neorv32_top.vhd:1031:38  */
  assign n769_o = io_acc & n768_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:1031:70  */
  assign n770_o = p_bus[99:96];
  /* ../neorv32/rtl/core/neorv32_top.vhd:1031:74  */
  assign n772_o = n770_o == 4'b1111;
  /* ../neorv32/rtl/core/neorv32_top.vhd:1031:59  */
  assign n773_o = n769_o & n772_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:1031:18  */
  assign n774_o = n773_o ? 1'b1 : 1'b0;
  /* ../neorv32/rtl/core/neorv32_top.vhd:1196:23  */
  assign n785_o = p_bus[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:1199:23  */
  assign n786_o = p_bus[95:64];
  /* ../neorv32/rtl/core/neorv32_top.vhd:1200:17  */
  assign neorv32_mtime_inst_true_neorv32_mtime_inst_n787 = neorv32_mtime_inst_true_neorv32_mtime_inst_data_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:1201:17  */
  assign neorv32_mtime_inst_true_neorv32_mtime_inst_n788 = neorv32_mtime_inst_true_neorv32_mtime_inst_ack_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:1203:17  */
  assign neorv32_mtime_inst_true_neorv32_mtime_inst_n789 = neorv32_mtime_inst_true_neorv32_mtime_inst_irq_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:1191:5  */
  neorv32_mtime neorv32_mtime_inst_true_neorv32_mtime_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_int),
    .addr_i(n785_o),
    .rden_i(io_rden),
    .wren_i(io_wren),
    .data_i(n786_o),
    .data_o(neorv32_mtime_inst_true_neorv32_mtime_inst_data_o),
    .ack_o(neorv32_mtime_inst_true_neorv32_mtime_inst_ack_o),
    .irq_o(neorv32_mtime_inst_true_neorv32_mtime_inst_irq_o));
  /* ../neorv32/rtl/core/neorv32_top.vhd:1230:28  */
  assign n797_o = p_bus[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:1233:28  */
  assign n798_o = p_bus[95:64];
  /* ../neorv32/rtl/core/neorv32_top.vhd:1234:22  */
  assign neorv32_uart0_inst_true_neorv32_uart0_inst_n799 = neorv32_uart0_inst_true_neorv32_uart0_inst_data_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:1235:22  */
  assign neorv32_uart0_inst_true_neorv32_uart0_inst_n800 = neorv32_uart0_inst_true_neorv32_uart0_inst_ack_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:1237:22  */
  assign neorv32_uart0_inst_true_neorv32_uart0_inst_n801 = neorv32_uart0_inst_true_neorv32_uart0_inst_clkgen_en_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:1240:22  */
  assign neorv32_uart0_inst_true_neorv32_uart0_inst_n802 = neorv32_uart0_inst_true_neorv32_uart0_inst_uart_txd_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:1243:22  */
  assign neorv32_uart0_inst_true_neorv32_uart0_inst_n803 = neorv32_uart0_inst_true_neorv32_uart0_inst_uart_rts_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:1246:22  */
  assign neorv32_uart0_inst_true_neorv32_uart0_inst_n804 = neorv32_uart0_inst_true_neorv32_uart0_inst_irq_rx_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:1247:22  */
  assign neorv32_uart0_inst_true_neorv32_uart0_inst_n805 = neorv32_uart0_inst_true_neorv32_uart0_inst_irq_tx_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:1220:5  */
  neorv32_uart_256_256_bf8b4530d8d246dd74ac53a13471bba17941dff7 neorv32_uart0_inst_true_neorv32_uart0_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_int),
    .addr_i(n797_o),
    .rden_i(io_rden),
    .wren_i(io_wren),
    .data_i(n798_o),
    .clkgen_i(clk_gen),
    .uart_rxd_i(uart0_rxd_i),
    .uart_cts_i(uart0_cts_i),
    .data_o(neorv32_uart0_inst_true_neorv32_uart0_inst_data_o),
    .ack_o(neorv32_uart0_inst_true_neorv32_uart0_inst_ack_o),
    .clkgen_en_o(neorv32_uart0_inst_true_neorv32_uart0_inst_clkgen_en_o),
    .uart_txd_o(neorv32_uart0_inst_true_neorv32_uart0_inst_uart_txd_o),
    .uart_rts_o(neorv32_uart0_inst_true_neorv32_uart0_inst_uart_rts_o),
    .irq_rx_o(neorv32_uart0_inst_true_neorv32_uart0_inst_irq_rx_o),
    .irq_tx_o(neorv32_uart0_inst_true_neorv32_uart0_inst_irq_tx_o));
  /* ../neorv32/rtl/core/neorv32_top.vhd:1656:21  */
  assign n846_o = p_bus[31:0];
  /* ../neorv32/rtl/core/neorv32_top.vhd:1659:15  */
  assign neorv32_sysinfo_inst_n847 = neorv32_sysinfo_inst_data_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:1660:15  */
  assign neorv32_sysinfo_inst_n848 = neorv32_sysinfo_inst_ack_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:1661:15  */
  assign neorv32_sysinfo_inst_n849 = neorv32_sysinfo_inst_err_o; // (signal)
  /* ../neorv32/rtl/core/neorv32_top.vhd:1607:3  */
  neorv32_sysinfo_5000000_0_1024_2048_4_64_1_4_64_0_0_0_c00c06f0c8f7e7aa711090f9c2d219a9079d700c neorv32_sysinfo_inst (
    .clk_i(clk_i),
    .addr_i(n846_o),
    .rden_i(io_rden),
    .wren_i(io_wren),
    .data_o(neorv32_sysinfo_inst_data_o),
    .ack_o(neorv32_sysinfo_inst_ack_o),
    .err_o(neorv32_sysinfo_inst_err_o));
  /* ../neorv32/rtl/core/neorv32_top.vhd:449:5  */
  always @(negedge clk_i or posedge n145_o)
    if (n145_o)
      n859_q <= 4'b0000;
    else
      n859_q <= n157_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:449:5  */
  always @(negedge clk_i or posedge n145_o)
    if (n145_o)
      n861_q <= 1'b0;
    else
      n861_q <= n189_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:473:5  */
  always @(posedge clk_i or posedge n204_o)
    if (n204_o)
      n862_q <= 12'b000000000000;
    else
      n862_q <= n239_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:473:5  */
  always @(posedge clk_i or posedge n204_o)
    if (n204_o)
      n863_q <= 12'b000000000000;
    else
      n863_q <= clk_div;
  /* ../neorv32/rtl/core/neorv32_top.vhd:469:5  */
  assign n864_o = {n281_o, n277_o, n273_o, n269_o, n265_o, n261_o, n257_o, n253_o};
  /* ../neorv32/rtl/core/neorv32_top.vhd:469:5  */
  assign n865_o = {onewire_cg_en, xip_cg_en, gptmr_cg_en, neoled_cg_en, cfs_cg_en, pwm_cg_en, twi_cg_en, spi_cg_en, uart1_cg_en, uart0_cg_en, wdt_cg_en};
  /* ../neorv32/rtl/core/neorv32_top.vhd:473:5  */
  always @(posedge clk_i or posedge n204_o)
    if (n204_o)
      n866_q <= 1'b0;
    else
      n866_q <= n235_o;
  /* ../neorv32/rtl/core/neorv32_top.vhd:444:5  */
  assign n868_o = {neorv32_cpu_inst_n290, 1'b0, 1'b1, neorv32_cpu_inst_n289, n341_o, n340_o, neorv32_cpu_inst_n286, n338_o, neorv32_cpu_inst_n284};
  /* ../neorv32/rtl/core/neorv32_top.vhd:444:5  */
  assign n869_o = {n342_o, 1'b0, 1'b0, 1'b0, neorv32_busswitch_inst_n376, neorv32_busswitch_inst_n375, n339_o, neorv32_busswitch_inst_n370, n337_o};
  /* ../neorv32/rtl/core/neorv32_top.vhd:444:5  */
  assign n870_o = {neorv32_cpu_inst_n300, 1'b0, 1'b0, neorv32_cpu_inst_n299, n353_o, n352_o, neorv32_cpu_inst_n296, neorv32_cpu_inst_n295, neorv32_cpu_inst_n294, neorv32_cpu_inst_n293, n347_o, neorv32_cpu_inst_n291};
  /* ../neorv32/rtl/core/neorv32_top.vhd:444:5  */
  assign n871_o = {n354_o, 1'b0, 1'b0, 1'b0, neorv32_busswitch_inst_n366, neorv32_busswitch_inst_n365, n351_o, n350_o, n349_o, n348_o, neorv32_busswitch_inst_n360, n346_o};
  assign n872_o = {neorv32_busswitch_inst_n377, neorv32_busswitch_inst_n378, neorv32_busswitch_inst_n379, n417_o, n643_o, n640_o, neorv32_busswitch_inst_n385, neorv32_busswitch_inst_n384, neorv32_busswitch_inst_n383, neorv32_busswitch_inst_n382, n637_o, neorv32_busswitch_inst_n380};
  assign n874_o = {1'b0, neorv32_bus_keeper_inst_n648, neorv32_bus_keeper_inst_n647, neorv32_int_imem_inst_true_neorv32_int_imem_inst_n669, neorv32_int_imem_inst_true_neorv32_int_imem_inst_n668, neorv32_int_imem_inst_true_neorv32_int_imem_inst_n667, 1'b0, neorv32_int_dmem_inst_true_neorv32_int_dmem_inst_n682, neorv32_int_dmem_inst_true_neorv32_int_dmem_inst_n681, neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_n693, neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_n692, neorv32_boot_rom_inst_true_neorv32_boot_rom_inst_n691, neorv32_wishbone_inst_true_neorv32_wishbone_inst_n708, neorv32_wishbone_inst_true_neorv32_wishbone_inst_n707, neorv32_wishbone_inst_true_neorv32_wishbone_inst_n706, 34'b0000000000000000000000000000000000, 1'b0, neorv32_mtime_inst_true_neorv32_mtime_inst_n788, neorv32_mtime_inst_true_neorv32_mtime_inst_n787, 1'b0, neorv32_uart0_inst_true_neorv32_uart0_inst_n800, neorv32_uart0_inst_true_neorv32_uart0_inst_n799, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, neorv32_sysinfo_inst_n849, neorv32_sysinfo_inst_n848, neorv32_sysinfo_inst_n847, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000};
  assign n875_o = {1'b0, 1'b0, onewire_irq, gptmr_irq, sdi_irq, 1'b0, neoled_irq, xirq_irq, twi_irq, spi_irq, uart1_tx_irq, uart1_rx_irq, uart0_tx_irq, uart0_rx_irq, cfs_irq, wdt_irq};
endmodule

module neorv32_verilog_wrapper
  (input  clk_i,
   input  rstn_i,
   input  uart0_rxd_i,
   input  [31:0] wb_dat_i,
   input  wb_ack_i,
   output uart0_txd_o,
   output [31:0] wb_adr_o,
   output [31:0] wb_dat_o,
   output wb_we_o,
   output [3:0] wb_sel_o,
   output wb_stb_o,
   output wb_cyc_o);
  localparam n7_o = 1'bX;
  localparam n8_o = 1'bX;
  localparam n9_o = 1'bX;
  localparam n11_o = 1'bX;
  wire [31:0] neorv32_top_inst_n13;
  wire [31:0] neorv32_top_inst_n14;
  wire neorv32_top_inst_n15;
  wire [3:0] neorv32_top_inst_n16;
  wire neorv32_top_inst_n17;
  wire neorv32_top_inst_n18;
  localparam n19_o = 1'b0;
  localparam n24_o = 1'b0;
  localparam [63:0] n27_o = 64'bX;
  wire neorv32_top_inst_n28;
  localparam n30_o = 1'b0;
  localparam n32_o = 1'bX;
  localparam n34_o = 1'b0;
  localparam n37_o = 1'bX;
  localparam n39_o = 1'bX;
  localparam n41_o = 1'bX;
  localparam n42_o = 1'b1;
  localparam n43_o = 1'b1;
  localparam n45_o = 1'b1;
  localparam n47_o = 1'b1;
  localparam [31:0] n50_o = 32'bX;
  localparam [31:0] n53_o = 32'b00000000000000000000000000000000;
  localparam n54_o = 1'b0;
  localparam n55_o = 1'b0;
  localparam n56_o = 1'b0;
  wire neorv32_top_inst_jtag_tdo_o;
  wire [2:0] neorv32_top_inst_wb_tag_o;
  wire [31:0] neorv32_top_inst_wb_adr_o;
  wire [31:0] neorv32_top_inst_wb_dat_o;
  wire neorv32_top_inst_wb_we_o;
  wire [3:0] neorv32_top_inst_wb_sel_o;
  wire neorv32_top_inst_wb_stb_o;
  wire neorv32_top_inst_wb_cyc_o;
  wire neorv32_top_inst_fence_o;
  wire neorv32_top_inst_fencei_o;
  wire neorv32_top_inst_xip_csn_o;
  wire neorv32_top_inst_xip_clk_o;
  wire neorv32_top_inst_xip_dat_o;
  wire [63:0] neorv32_top_inst_gpio_o;
  wire neorv32_top_inst_uart0_txd_o;
  wire neorv32_top_inst_uart0_rts_o;
  wire neorv32_top_inst_uart1_txd_o;
  wire neorv32_top_inst_uart1_rts_o;
  wire neorv32_top_inst_spi_clk_o;
  wire neorv32_top_inst_spi_dat_o;
  wire [7:0] neorv32_top_inst_spi_csn_o;
  wire neorv32_top_inst_sdi_dat_o;
  wire neorv32_top_inst_twi_sda_o;
  wire neorv32_top_inst_twi_scl_o;
  wire neorv32_top_inst_onewire_o;
  wire [11:0] neorv32_top_inst_pwm_o;
  wire [31:0] neorv32_top_inst_cfs_out_o;
  wire neorv32_top_inst_neoled_o;
  assign uart0_txd_o = neorv32_top_inst_n28;
  assign wb_adr_o = neorv32_top_inst_n13;
  assign wb_dat_o = neorv32_top_inst_n14;
  assign wb_we_o = neorv32_top_inst_n15;
  assign wb_sel_o = neorv32_top_inst_n16;
  assign wb_stb_o = neorv32_top_inst_n17;
  assign wb_cyc_o = neorv32_top_inst_n18;
  /* ./neorv32_verilog_wrapper.vhd:63:20  */
  assign neorv32_top_inst_n13 = neorv32_top_inst_wb_adr_o; // (signal)
  /* ./neorv32_verilog_wrapper.vhd:65:20  */
  assign neorv32_top_inst_n14 = neorv32_top_inst_wb_dat_o; // (signal)
  /* ./neorv32_verilog_wrapper.vhd:66:20  */
  assign neorv32_top_inst_n15 = neorv32_top_inst_wb_we_o; // (signal)
  /* ./neorv32_verilog_wrapper.vhd:67:20  */
  assign neorv32_top_inst_n16 = neorv32_top_inst_wb_sel_o; // (signal)
  /* ./neorv32_verilog_wrapper.vhd:68:20  */
  assign neorv32_top_inst_n17 = neorv32_top_inst_wb_stb_o; // (signal)
  /* ./neorv32_verilog_wrapper.vhd:69:20  */
  assign neorv32_top_inst_n18 = neorv32_top_inst_wb_cyc_o; // (signal)
  /* ./neorv32_verilog_wrapper.vhd:60:20  */
  assign neorv32_top_inst_n28 = neorv32_top_inst_uart0_txd_o; // (signal)
  /* ./neorv32_verilog_wrapper.vhd:31:3  */
  neorv32_top_5000000_1_0_4_0_40_1024_2048_4_64_1_4_64_255_0_0_256_256_1_1_1_0_0_1_32_32_1_69ad7886168de6916fb842204ba7129434750df3 neorv32_top_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .jtag_trst_i(n7_o),
    .jtag_tck_i(n8_o),
    .jtag_tdi_i(n9_o),
    .jtag_tms_i(n11_o),
    .wb_dat_i(wb_dat_i),
    .wb_ack_i(wb_ack_i),
    .wb_err_i(n19_o),
    .xip_dat_i(n24_o),
    .gpio_i(n27_o),
    .uart0_rxd_i(uart0_rxd_i),
    .uart0_cts_i(n30_o),
    .uart1_rxd_i(n32_o),
    .uart1_cts_i(n34_o),
    .spi_dat_i(n37_o),
    .sdi_clk_i(n39_o),
    .sdi_dat_i(n41_o),
    .sdi_csn_i(n42_o),
    .twi_sda_i(n43_o),
    .twi_scl_i(n45_o),
    .onewire_i(n47_o),
    .cfs_in_i(n50_o),
    .xirq_i(n53_o),
    .mtime_irq_i(n54_o),
    .msw_irq_i(n55_o),
    .mext_irq_i(n56_o),
    .jtag_tdo_o(),
    .wb_tag_o(),
    .wb_adr_o(neorv32_top_inst_wb_adr_o),
    .wb_dat_o(neorv32_top_inst_wb_dat_o),
    .wb_we_o(neorv32_top_inst_wb_we_o),
    .wb_sel_o(neorv32_top_inst_wb_sel_o),
    .wb_stb_o(neorv32_top_inst_wb_stb_o),
    .wb_cyc_o(neorv32_top_inst_wb_cyc_o),
    .fence_o(),
    .fencei_o(),
    .xip_csn_o(),
    .xip_clk_o(),
    .xip_dat_o(),
    .gpio_o(),
    .uart0_txd_o(neorv32_top_inst_uart0_txd_o),
    .uart0_rts_o(),
    .uart1_txd_o(),
    .uart1_rts_o(),
    .spi_clk_o(),
    .spi_dat_o(),
    .spi_csn_o(),
    .sdi_dat_o(),
    .twi_sda_o(),
    .twi_scl_o(),
    .onewire_o(),
    .pwm_o(),
    .cfs_out_o(),
    .neoled_o());
endmodule

